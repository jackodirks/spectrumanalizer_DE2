---------------------------------------------------------------------------------------------------
--- State Machine Template ------------------------------------------------------------------------
---------------------------------------------------------------------------------------------------
-- Author  : PelJH          
-- Date    : 15-09-2010     
-- Version : V1.0
-- Name    : statemachine.vhd
---------------------------------------------------------------------------------------------------
-- Description:             
-- This template is meant to be used by students of the HWP01 course at the Hogeschool Rotterdam
-- It implements a basic FSM in VHDL. Please note that there are many other ways to do this.
-- Students may also use the FSM templates by Altera that can be found in the template library of
-- Quartus. Also other templates are allowed that can be found in books and online. It is mandatory,
-- however, that the FSM templates used give a good vice-versa overview in relation to the FSM 
-- diagram that must be drawn for the assignments.
---------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ADC_sampler is 
	port	( 	
				-- clock and reset
				CLOCK_50:  	in std_logic;
				CLOCK_27:	IN STD_LOGIC;
				reset: 		in std_logic;
				
				-- list of inputs
				CONTROL:   	in std_logic;								--start/stop input
				--KEY:   		in std_logic_vector(0 downto 0);
				ADC_BUSY:	in std_logic;
				ADC:    		inout std_logic_vector(11 downto 0);
				
				-- list of outputs
				DONE:    	out std_logic;								--samples are ready
				--LEDR:   		out std_logic_vector(7 downto 0);
				LEDG:   		out std_logic_vector(7 downto 0);
				ADC_CLKIN:  out std_logic;	
				ADC_CONVST: out std_logic;
				ADC_WB: 		out std_logic;
				ADC_WR:		out std_logic;
				ADC_RD: 		out std_logic;
				ADC_CS: 		out std_logic;	
				
				samples:   out std_logic_vector(20479 DOWNTO 0)
			);
end ADC_sampler;

architecture ADC_sampler of ADC_sampler is

component ADC_CLK_prescaler IS
	PORT
	(
		areset		: IN STD_LOGIC  := '0';
		inclk0		: IN STD_LOGIC  := '0';
		c0			: OUT STD_LOGIC ;
		locked		: OUT STD_LOGIC 
	);
END component;

component ADC_setup_timer IS
	PORT
	(
		clock_50m	: IN STD_LOGIC;
		reset		: IN STD_LOGIC;
		done		: OUT STD_LOGIC
	);
END component;

component ADC_sample_timer IS
	PORT
	(
		clock_50m: IN STD_LOGIC;
		reset		: IN STD_LOGIC;
		done		: OUT STD_LOGIC
	);
END component;

component ADC_sample_counter IS
	PORT
	(
		clock_50m	: IN STD_LOGIC;
		increment	: IN STD_LOGIC;
		reset		: IN STD_LOGIC;
		done		: OUT STD_LOGIC;
		count		: OUT STD_LOGIC_VECTOR(11 downto 0)
	);
END component;

signal CLOCK_10	: STD_LOGIC;
SIGNAL timer_reset: STD_LOGIC ;
SIGNAL timer_done	: STD_LOGIC ;

SIGNAL setup_timer_reset: STD_LOGIC ;
SIGNAL setup_timer_done	: STD_LOGIC ;

SIGNAL sample_counter_increment : STD_LOGIC ;
SIGNAL sample_counter_reset: STD_LOGIC ;
SIGNAL sample_counter_done	: STD_LOGIC ;
Signal sample_count : STD_LOGIC_VECTOR(11 downto 0);


-------------------------------------------------------------------
-- state definitions and signals ----------------------------------
-------------------------------------------------------------------
	type state is ( state_0,
					state_1,
					state_2,
					state_3,
					state_4,
					state_5);
						
	signal present_state, next_state: state;
	attribute enum_encoding : string;
	attribute enum_encoding of state : type is "gray";

begin

	ADC_CLKIN	<= CLOCK_10;

	prescaler : ADC_CLK_prescaler
	port map
	(
		inclk0 => CLOCK_27, 
		c0 => CLOCK_10
	);

	timer : ADC_sample_timer
	port map
	(
		clock_50m => CLOCK_50,
		reset	=> timer_reset,
		done => timer_done
	);
	
	setup_timer : ADC_setup_timer
	port map
	(
		clock_50m => CLOCK_50,
		reset	=> setup_timer_reset,
		done => setup_timer_done
	);
	
	sample_counter : ADC_sample_counter
	port map
	(
		clock_50m => CLOCK_50,
		increment => sample_counter_increment,
		reset	=> sample_counter_reset,
		done => sample_counter_done,
		count => sample_count
	);

-------------------------------------------------------------------
-- sequential part of the statemachine ----------------------------
-------------------------------------------------------------------
	process(reset, CLOCK_50)
	begin
		if (reset = '0') 
		then
			present_state <= state_0;
		elsif (rising_edge(CLOCK_50)) 
		then
			present_state <= next_state;
		end if;
	end process;
-------------------------------------------------------------------
	
-------------------------------------------------------------------
-- combinatorial part of the statemachine -------------------------
-------------------------------------------------------------------
	process (--KEY,
				ADC,
				-- add other inputs to use for next state testing 
				-- or to generate outputs with
				present_state,
				timer_done,
				setup_timer_done,
				sample_counter_done,
				sample_count,
				CONTROL
				)
				
	------------------------------- gen by c
	variable temp: std_logic_vector(20479 downto 0) := (OTHERS => '0');
	----------------------------------------
	begin
	
-- Default values of outputs
			DONE			<= '0';
			ADC_CONVST	<= '0';
			ADC_WB		<= '1';
			ADC_WR		<= '1';
			ADC_RD		<= '1';
			ADC_CS		<= '1';
			LEDG 			<= "00000000";
			ADC 			<= "ZZZZZZZZZZZZ";
			timer_reset <= '1';
			setup_timer_reset <= '1';
			
			sample_counter_increment <= '0';
			sample_counter_reset <= '1';
		
				ADC 			<= "ZZZZZZZZZZZZ";
			--LEDR(7 downto 0) <= "00000000";
		
		case present_state is
--------------------------------------
-- state 0  INIT                    --
--------------------------------------
			when state_0 =>
				--------------------------
				-- determine next state --
				--------------------------
				if (setup_timer_done = '1')
				then
					next_state <= state_1;
				else
					next_state <= present_state;
				end if;
				--------------------------
				--  determine outputs   --
				--------------------------
				DONE			<= '0';
				ADC_CONVST	<= '1';
				ADC_WB		<= '1';
				ADC_WR		<= '0';
				ADC_RD		<= '1';
				ADC_CS		<= '0';
				LEDG 			<= "00000001";
				ADC 			<= "000000010110"; -- tows compliment <= "001000010110";
				timer_reset <= '1';
				setup_timer_reset <= '0';	
							
				sample_counter_increment <= '0';
				sample_counter_reset <= '1';
		
--------------------------------------
-- state 1  IDLE                    --
--------------------------------------
			when state_1 =>
				--------------------------
				-- determine next state --
				--------------------------
				if (CONTROL = '1') --START
				then
					next_state <= state_2;
				else
					next_state <= present_state;
				end if;
				--------------------------
				--  determine outputs   --
				--------------------------
				DONE			<= '0';
				ADC_CONVST	<= '1';
				ADC_WB		<= '1';
				ADC_WR		<= '1';
				ADC_RD		<= '1';
				ADC_CS		<= '0';
				ADC 			<= "ZZZZZZZZZZZZ";
				LEDG 			<= "00000010";
				timer_reset <= '1';
				setup_timer_reset <= '1';
							
				sample_counter_increment <= '0';
				sample_counter_reset <= '1';

--------------------------------------
-- state 2 sample wait              --
--------------------------------------
			when state_2 =>
				--------------------------
				-- determine next state --
				--------------------------
				if (timer_done = '1')
				then
					next_state <= state_3;
				else
					next_state <= present_state;
				end if;
				--------------------------
				--  determine outputs   --
				--------------------------
				DONE			<= '0';
				ADC_CONVST	<= '0';
				ADC_WB		<= '1';
				ADC_WR		<= '1';
				ADC_RD		<= '0';
				ADC_CS		<= '0';
				ADC 			<= "ZZZZZZZZZZZZ";
				LEDG 			<= "00000100";
				timer_reset <= '0';
				setup_timer_reset <= '1';
				
				sample_counter_increment <= '0';
				sample_counter_reset <= '0';
--------------------------------------
-- state 3 grab sample              --
--------------------------------------
			when state_3 =>
				--------------------------
				-- determine next state --
				--------------------------
				if (timer_done = '0') then
					if (sample_counter_done = '0') then
						next_state <= state_4;
					else
						next_state <= state_5;
					end if;
				else
					next_state <= present_state;
				ADC 			<= "ZZZZZZZZZZZZ";
				end if;
				--------------------------
				--  determine outputs   --
				--------------------------
				DONE			<= '0';
				ADC_CONVST	<= '1';
				ADC_WB		<= '1';
				ADC_WR		<= '1';
				ADC_RD		<= '0';
				ADC_CS		<= '0';
				ADC 			<= "ZZZZZZZZZZZZ";
				--LEDG 			<= "00001000";
				timer_reset <= '1';
				setup_timer_reset <= '1';
				
				sample_counter_increment <= '0';
				sample_counter_reset <= '0';
				--TEMP
				LEDG <= ADC(11 DOWNTO 4);
				
				case to_integer(unsigned(sample_count)) is
					------------------------------- gen by c	
					when 0 => temp(9 downto 0) := ADC(11 downto 2);
					when 1 => temp(19 downto 10) := ADC(11 downto 2);
					when 2 => temp(29 downto 20) := ADC(11 downto 2);
					when 3 => temp(39 downto 30) := ADC(11 downto 2);
					when 4 => temp(49 downto 40) := ADC(11 downto 2);
					when 5 => temp(59 downto 50) := ADC(11 downto 2);
					when 6 => temp(69 downto 60) := ADC(11 downto 2);
					when 7 => temp(79 downto 70) := ADC(11 downto 2);
					when 8 => temp(89 downto 80) := ADC(11 downto 2);
					when 9 => temp(99 downto 90) := ADC(11 downto 2);
					when 10 => temp(109 downto 100) := ADC(11 downto 2);
					when 11 => temp(119 downto 110) := ADC(11 downto 2);
					when 12 => temp(129 downto 120) := ADC(11 downto 2);
					when 13 => temp(139 downto 130) := ADC(11 downto 2);
					when 14 => temp(149 downto 140) := ADC(11 downto 2);
					when 15 => temp(159 downto 150) := ADC(11 downto 2);
					when 16 => temp(169 downto 160) := ADC(11 downto 2);
					when 17 => temp(179 downto 170) := ADC(11 downto 2);
					when 18 => temp(189 downto 180) := ADC(11 downto 2);
					when 19 => temp(199 downto 190) := ADC(11 downto 2);
					when 20 => temp(209 downto 200) := ADC(11 downto 2);
					when 21 => temp(219 downto 210) := ADC(11 downto 2);
					when 22 => temp(229 downto 220) := ADC(11 downto 2);
					when 23 => temp(239 downto 230) := ADC(11 downto 2);
					when 24 => temp(249 downto 240) := ADC(11 downto 2);
					when 25 => temp(259 downto 250) := ADC(11 downto 2);
					when 26 => temp(269 downto 260) := ADC(11 downto 2);
					when 27 => temp(279 downto 270) := ADC(11 downto 2);
					when 28 => temp(289 downto 280) := ADC(11 downto 2);
					when 29 => temp(299 downto 290) := ADC(11 downto 2);
					when 30 => temp(309 downto 300) := ADC(11 downto 2);
					when 31 => temp(319 downto 310) := ADC(11 downto 2);
					when 32 => temp(329 downto 320) := ADC(11 downto 2);
					when 33 => temp(339 downto 330) := ADC(11 downto 2);
					when 34 => temp(349 downto 340) := ADC(11 downto 2);
					when 35 => temp(359 downto 350) := ADC(11 downto 2);
					when 36 => temp(369 downto 360) := ADC(11 downto 2);
					when 37 => temp(379 downto 370) := ADC(11 downto 2);
					when 38 => temp(389 downto 380) := ADC(11 downto 2);
					when 39 => temp(399 downto 390) := ADC(11 downto 2);
					when 40 => temp(409 downto 400) := ADC(11 downto 2);
					when 41 => temp(419 downto 410) := ADC(11 downto 2);
					when 42 => temp(429 downto 420) := ADC(11 downto 2);
					when 43 => temp(439 downto 430) := ADC(11 downto 2);
					when 44 => temp(449 downto 440) := ADC(11 downto 2);
					when 45 => temp(459 downto 450) := ADC(11 downto 2);
					when 46 => temp(469 downto 460) := ADC(11 downto 2);
					when 47 => temp(479 downto 470) := ADC(11 downto 2);
					when 48 => temp(489 downto 480) := ADC(11 downto 2);
					when 49 => temp(499 downto 490) := ADC(11 downto 2);
					when 50 => temp(509 downto 500) := ADC(11 downto 2);
					when 51 => temp(519 downto 510) := ADC(11 downto 2);
					when 52 => temp(529 downto 520) := ADC(11 downto 2);
					when 53 => temp(539 downto 530) := ADC(11 downto 2);
					when 54 => temp(549 downto 540) := ADC(11 downto 2);
					when 55 => temp(559 downto 550) := ADC(11 downto 2);
					when 56 => temp(569 downto 560) := ADC(11 downto 2);
					when 57 => temp(579 downto 570) := ADC(11 downto 2);
					when 58 => temp(589 downto 580) := ADC(11 downto 2);
					when 59 => temp(599 downto 590) := ADC(11 downto 2);
					when 60 => temp(609 downto 600) := ADC(11 downto 2);
					when 61 => temp(619 downto 610) := ADC(11 downto 2);
					when 62 => temp(629 downto 620) := ADC(11 downto 2);
					when 63 => temp(639 downto 630) := ADC(11 downto 2);
					when 64 => temp(649 downto 640) := ADC(11 downto 2);
					when 65 => temp(659 downto 650) := ADC(11 downto 2);
					when 66 => temp(669 downto 660) := ADC(11 downto 2);
					when 67 => temp(679 downto 670) := ADC(11 downto 2);
					when 68 => temp(689 downto 680) := ADC(11 downto 2);
					when 69 => temp(699 downto 690) := ADC(11 downto 2);
					when 70 => temp(709 downto 700) := ADC(11 downto 2);
					when 71 => temp(719 downto 710) := ADC(11 downto 2);
					when 72 => temp(729 downto 720) := ADC(11 downto 2);
					when 73 => temp(739 downto 730) := ADC(11 downto 2);
					when 74 => temp(749 downto 740) := ADC(11 downto 2);
					when 75 => temp(759 downto 750) := ADC(11 downto 2);
					when 76 => temp(769 downto 760) := ADC(11 downto 2);
					when 77 => temp(779 downto 770) := ADC(11 downto 2);
					when 78 => temp(789 downto 780) := ADC(11 downto 2);
					when 79 => temp(799 downto 790) := ADC(11 downto 2);
					when 80 => temp(809 downto 800) := ADC(11 downto 2);
					when 81 => temp(819 downto 810) := ADC(11 downto 2);
					when 82 => temp(829 downto 820) := ADC(11 downto 2);
					when 83 => temp(839 downto 830) := ADC(11 downto 2);
					when 84 => temp(849 downto 840) := ADC(11 downto 2);
					when 85 => temp(859 downto 850) := ADC(11 downto 2);
					when 86 => temp(869 downto 860) := ADC(11 downto 2);
					when 87 => temp(879 downto 870) := ADC(11 downto 2);
					when 88 => temp(889 downto 880) := ADC(11 downto 2);
					when 89 => temp(899 downto 890) := ADC(11 downto 2);
					when 90 => temp(909 downto 900) := ADC(11 downto 2);
					when 91 => temp(919 downto 910) := ADC(11 downto 2);
					when 92 => temp(929 downto 920) := ADC(11 downto 2);
					when 93 => temp(939 downto 930) := ADC(11 downto 2);
					when 94 => temp(949 downto 940) := ADC(11 downto 2);
					when 95 => temp(959 downto 950) := ADC(11 downto 2);
					when 96 => temp(969 downto 960) := ADC(11 downto 2);
					when 97 => temp(979 downto 970) := ADC(11 downto 2);
					when 98 => temp(989 downto 980) := ADC(11 downto 2);
					when 99 => temp(999 downto 990) := ADC(11 downto 2);
					when 100 => temp(1009 downto 1000) := ADC(11 downto 2);
					when 101 => temp(1019 downto 1010) := ADC(11 downto 2);
					when 102 => temp(1029 downto 1020) := ADC(11 downto 2);
					when 103 => temp(1039 downto 1030) := ADC(11 downto 2);
					when 104 => temp(1049 downto 1040) := ADC(11 downto 2);
					when 105 => temp(1059 downto 1050) := ADC(11 downto 2);
					when 106 => temp(1069 downto 1060) := ADC(11 downto 2);
					when 107 => temp(1079 downto 1070) := ADC(11 downto 2);
					when 108 => temp(1089 downto 1080) := ADC(11 downto 2);
					when 109 => temp(1099 downto 1090) := ADC(11 downto 2);
					when 110 => temp(1109 downto 1100) := ADC(11 downto 2);
					when 111 => temp(1119 downto 1110) := ADC(11 downto 2);
					when 112 => temp(1129 downto 1120) := ADC(11 downto 2);
					when 113 => temp(1139 downto 1130) := ADC(11 downto 2);
					when 114 => temp(1149 downto 1140) := ADC(11 downto 2);
					when 115 => temp(1159 downto 1150) := ADC(11 downto 2);
					when 116 => temp(1169 downto 1160) := ADC(11 downto 2);
					when 117 => temp(1179 downto 1170) := ADC(11 downto 2);
					when 118 => temp(1189 downto 1180) := ADC(11 downto 2);
					when 119 => temp(1199 downto 1190) := ADC(11 downto 2);
					when 120 => temp(1209 downto 1200) := ADC(11 downto 2);
					when 121 => temp(1219 downto 1210) := ADC(11 downto 2);
					when 122 => temp(1229 downto 1220) := ADC(11 downto 2);
					when 123 => temp(1239 downto 1230) := ADC(11 downto 2);
					when 124 => temp(1249 downto 1240) := ADC(11 downto 2);
					when 125 => temp(1259 downto 1250) := ADC(11 downto 2);
					when 126 => temp(1269 downto 1260) := ADC(11 downto 2);
					when 127 => temp(1279 downto 1270) := ADC(11 downto 2);
					when 128 => temp(1289 downto 1280) := ADC(11 downto 2);
					when 129 => temp(1299 downto 1290) := ADC(11 downto 2);
					when 130 => temp(1309 downto 1300) := ADC(11 downto 2);
					when 131 => temp(1319 downto 1310) := ADC(11 downto 2);
					when 132 => temp(1329 downto 1320) := ADC(11 downto 2);
					when 133 => temp(1339 downto 1330) := ADC(11 downto 2);
					when 134 => temp(1349 downto 1340) := ADC(11 downto 2);
					when 135 => temp(1359 downto 1350) := ADC(11 downto 2);
					when 136 => temp(1369 downto 1360) := ADC(11 downto 2);
					when 137 => temp(1379 downto 1370) := ADC(11 downto 2);
					when 138 => temp(1389 downto 1380) := ADC(11 downto 2);
					when 139 => temp(1399 downto 1390) := ADC(11 downto 2);
					when 140 => temp(1409 downto 1400) := ADC(11 downto 2);
					when 141 => temp(1419 downto 1410) := ADC(11 downto 2);
					when 142 => temp(1429 downto 1420) := ADC(11 downto 2);
					when 143 => temp(1439 downto 1430) := ADC(11 downto 2);
					when 144 => temp(1449 downto 1440) := ADC(11 downto 2);
					when 145 => temp(1459 downto 1450) := ADC(11 downto 2);
					when 146 => temp(1469 downto 1460) := ADC(11 downto 2);
					when 147 => temp(1479 downto 1470) := ADC(11 downto 2);
					when 148 => temp(1489 downto 1480) := ADC(11 downto 2);
					when 149 => temp(1499 downto 1490) := ADC(11 downto 2);
					when 150 => temp(1509 downto 1500) := ADC(11 downto 2);
					when 151 => temp(1519 downto 1510) := ADC(11 downto 2);
					when 152 => temp(1529 downto 1520) := ADC(11 downto 2);
					when 153 => temp(1539 downto 1530) := ADC(11 downto 2);
					when 154 => temp(1549 downto 1540) := ADC(11 downto 2);
					when 155 => temp(1559 downto 1550) := ADC(11 downto 2);
					when 156 => temp(1569 downto 1560) := ADC(11 downto 2);
					when 157 => temp(1579 downto 1570) := ADC(11 downto 2);
					when 158 => temp(1589 downto 1580) := ADC(11 downto 2);
					when 159 => temp(1599 downto 1590) := ADC(11 downto 2);
					when 160 => temp(1609 downto 1600) := ADC(11 downto 2);
					when 161 => temp(1619 downto 1610) := ADC(11 downto 2);
					when 162 => temp(1629 downto 1620) := ADC(11 downto 2);
					when 163 => temp(1639 downto 1630) := ADC(11 downto 2);
					when 164 => temp(1649 downto 1640) := ADC(11 downto 2);
					when 165 => temp(1659 downto 1650) := ADC(11 downto 2);
					when 166 => temp(1669 downto 1660) := ADC(11 downto 2);
					when 167 => temp(1679 downto 1670) := ADC(11 downto 2);
					when 168 => temp(1689 downto 1680) := ADC(11 downto 2);
					when 169 => temp(1699 downto 1690) := ADC(11 downto 2);
					when 170 => temp(1709 downto 1700) := ADC(11 downto 2);
					when 171 => temp(1719 downto 1710) := ADC(11 downto 2);
					when 172 => temp(1729 downto 1720) := ADC(11 downto 2);
					when 173 => temp(1739 downto 1730) := ADC(11 downto 2);
					when 174 => temp(1749 downto 1740) := ADC(11 downto 2);
					when 175 => temp(1759 downto 1750) := ADC(11 downto 2);
					when 176 => temp(1769 downto 1760) := ADC(11 downto 2);
					when 177 => temp(1779 downto 1770) := ADC(11 downto 2);
					when 178 => temp(1789 downto 1780) := ADC(11 downto 2);
					when 179 => temp(1799 downto 1790) := ADC(11 downto 2);
					when 180 => temp(1809 downto 1800) := ADC(11 downto 2);
					when 181 => temp(1819 downto 1810) := ADC(11 downto 2);
					when 182 => temp(1829 downto 1820) := ADC(11 downto 2);
					when 183 => temp(1839 downto 1830) := ADC(11 downto 2);
					when 184 => temp(1849 downto 1840) := ADC(11 downto 2);
					when 185 => temp(1859 downto 1850) := ADC(11 downto 2);
					when 186 => temp(1869 downto 1860) := ADC(11 downto 2);
					when 187 => temp(1879 downto 1870) := ADC(11 downto 2);
					when 188 => temp(1889 downto 1880) := ADC(11 downto 2);
					when 189 => temp(1899 downto 1890) := ADC(11 downto 2);
					when 190 => temp(1909 downto 1900) := ADC(11 downto 2);
					when 191 => temp(1919 downto 1910) := ADC(11 downto 2);
					when 192 => temp(1929 downto 1920) := ADC(11 downto 2);
					when 193 => temp(1939 downto 1930) := ADC(11 downto 2);
					when 194 => temp(1949 downto 1940) := ADC(11 downto 2);
					when 195 => temp(1959 downto 1950) := ADC(11 downto 2);
					when 196 => temp(1969 downto 1960) := ADC(11 downto 2);
					when 197 => temp(1979 downto 1970) := ADC(11 downto 2);
					when 198 => temp(1989 downto 1980) := ADC(11 downto 2);
					when 199 => temp(1999 downto 1990) := ADC(11 downto 2);
					when 200 => temp(2009 downto 2000) := ADC(11 downto 2);
					when 201 => temp(2019 downto 2010) := ADC(11 downto 2);
					when 202 => temp(2029 downto 2020) := ADC(11 downto 2);
					when 203 => temp(2039 downto 2030) := ADC(11 downto 2);
					when 204 => temp(2049 downto 2040) := ADC(11 downto 2);
					when 205 => temp(2059 downto 2050) := ADC(11 downto 2);
					when 206 => temp(2069 downto 2060) := ADC(11 downto 2);
					when 207 => temp(2079 downto 2070) := ADC(11 downto 2);
					when 208 => temp(2089 downto 2080) := ADC(11 downto 2);
					when 209 => temp(2099 downto 2090) := ADC(11 downto 2);
					when 210 => temp(2109 downto 2100) := ADC(11 downto 2);
					when 211 => temp(2119 downto 2110) := ADC(11 downto 2);
					when 212 => temp(2129 downto 2120) := ADC(11 downto 2);
					when 213 => temp(2139 downto 2130) := ADC(11 downto 2);
					when 214 => temp(2149 downto 2140) := ADC(11 downto 2);
					when 215 => temp(2159 downto 2150) := ADC(11 downto 2);
					when 216 => temp(2169 downto 2160) := ADC(11 downto 2);
					when 217 => temp(2179 downto 2170) := ADC(11 downto 2);
					when 218 => temp(2189 downto 2180) := ADC(11 downto 2);
					when 219 => temp(2199 downto 2190) := ADC(11 downto 2);
					when 220 => temp(2209 downto 2200) := ADC(11 downto 2);
					when 221 => temp(2219 downto 2210) := ADC(11 downto 2);
					when 222 => temp(2229 downto 2220) := ADC(11 downto 2);
					when 223 => temp(2239 downto 2230) := ADC(11 downto 2);
					when 224 => temp(2249 downto 2240) := ADC(11 downto 2);
					when 225 => temp(2259 downto 2250) := ADC(11 downto 2);
					when 226 => temp(2269 downto 2260) := ADC(11 downto 2);
					when 227 => temp(2279 downto 2270) := ADC(11 downto 2);
					when 228 => temp(2289 downto 2280) := ADC(11 downto 2);
					when 229 => temp(2299 downto 2290) := ADC(11 downto 2);
					when 230 => temp(2309 downto 2300) := ADC(11 downto 2);
					when 231 => temp(2319 downto 2310) := ADC(11 downto 2);
					when 232 => temp(2329 downto 2320) := ADC(11 downto 2);
					when 233 => temp(2339 downto 2330) := ADC(11 downto 2);
					when 234 => temp(2349 downto 2340) := ADC(11 downto 2);
					when 235 => temp(2359 downto 2350) := ADC(11 downto 2);
					when 236 => temp(2369 downto 2360) := ADC(11 downto 2);
					when 237 => temp(2379 downto 2370) := ADC(11 downto 2);
					when 238 => temp(2389 downto 2380) := ADC(11 downto 2);
					when 239 => temp(2399 downto 2390) := ADC(11 downto 2);
					when 240 => temp(2409 downto 2400) := ADC(11 downto 2);
					when 241 => temp(2419 downto 2410) := ADC(11 downto 2);
					when 242 => temp(2429 downto 2420) := ADC(11 downto 2);
					when 243 => temp(2439 downto 2430) := ADC(11 downto 2);
					when 244 => temp(2449 downto 2440) := ADC(11 downto 2);
					when 245 => temp(2459 downto 2450) := ADC(11 downto 2);
					when 246 => temp(2469 downto 2460) := ADC(11 downto 2);
					when 247 => temp(2479 downto 2470) := ADC(11 downto 2);
					when 248 => temp(2489 downto 2480) := ADC(11 downto 2);
					when 249 => temp(2499 downto 2490) := ADC(11 downto 2);
					when 250 => temp(2509 downto 2500) := ADC(11 downto 2);
					when 251 => temp(2519 downto 2510) := ADC(11 downto 2);
					when 252 => temp(2529 downto 2520) := ADC(11 downto 2);
					when 253 => temp(2539 downto 2530) := ADC(11 downto 2);
					when 254 => temp(2549 downto 2540) := ADC(11 downto 2);
					when 255 => temp(2559 downto 2550) := ADC(11 downto 2);
					when 256 => temp(2569 downto 2560) := ADC(11 downto 2);
					when 257 => temp(2579 downto 2570) := ADC(11 downto 2);
					when 258 => temp(2589 downto 2580) := ADC(11 downto 2);
					when 259 => temp(2599 downto 2590) := ADC(11 downto 2);
					when 260 => temp(2609 downto 2600) := ADC(11 downto 2);
					when 261 => temp(2619 downto 2610) := ADC(11 downto 2);
					when 262 => temp(2629 downto 2620) := ADC(11 downto 2);
					when 263 => temp(2639 downto 2630) := ADC(11 downto 2);
					when 264 => temp(2649 downto 2640) := ADC(11 downto 2);
					when 265 => temp(2659 downto 2650) := ADC(11 downto 2);
					when 266 => temp(2669 downto 2660) := ADC(11 downto 2);
					when 267 => temp(2679 downto 2670) := ADC(11 downto 2);
					when 268 => temp(2689 downto 2680) := ADC(11 downto 2);
					when 269 => temp(2699 downto 2690) := ADC(11 downto 2);
					when 270 => temp(2709 downto 2700) := ADC(11 downto 2);
					when 271 => temp(2719 downto 2710) := ADC(11 downto 2);
					when 272 => temp(2729 downto 2720) := ADC(11 downto 2);
					when 273 => temp(2739 downto 2730) := ADC(11 downto 2);
					when 274 => temp(2749 downto 2740) := ADC(11 downto 2);
					when 275 => temp(2759 downto 2750) := ADC(11 downto 2);
					when 276 => temp(2769 downto 2760) := ADC(11 downto 2);
					when 277 => temp(2779 downto 2770) := ADC(11 downto 2);
					when 278 => temp(2789 downto 2780) := ADC(11 downto 2);
					when 279 => temp(2799 downto 2790) := ADC(11 downto 2);
					when 280 => temp(2809 downto 2800) := ADC(11 downto 2);
					when 281 => temp(2819 downto 2810) := ADC(11 downto 2);
					when 282 => temp(2829 downto 2820) := ADC(11 downto 2);
					when 283 => temp(2839 downto 2830) := ADC(11 downto 2);
					when 284 => temp(2849 downto 2840) := ADC(11 downto 2);
					when 285 => temp(2859 downto 2850) := ADC(11 downto 2);
					when 286 => temp(2869 downto 2860) := ADC(11 downto 2);
					when 287 => temp(2879 downto 2870) := ADC(11 downto 2);
					when 288 => temp(2889 downto 2880) := ADC(11 downto 2);
					when 289 => temp(2899 downto 2890) := ADC(11 downto 2);
					when 290 => temp(2909 downto 2900) := ADC(11 downto 2);
					when 291 => temp(2919 downto 2910) := ADC(11 downto 2);
					when 292 => temp(2929 downto 2920) := ADC(11 downto 2);
					when 293 => temp(2939 downto 2930) := ADC(11 downto 2);
					when 294 => temp(2949 downto 2940) := ADC(11 downto 2);
					when 295 => temp(2959 downto 2950) := ADC(11 downto 2);
					when 296 => temp(2969 downto 2960) := ADC(11 downto 2);
					when 297 => temp(2979 downto 2970) := ADC(11 downto 2);
					when 298 => temp(2989 downto 2980) := ADC(11 downto 2);
					when 299 => temp(2999 downto 2990) := ADC(11 downto 2);
					when 300 => temp(3009 downto 3000) := ADC(11 downto 2);
					when 301 => temp(3019 downto 3010) := ADC(11 downto 2);
					when 302 => temp(3029 downto 3020) := ADC(11 downto 2);
					when 303 => temp(3039 downto 3030) := ADC(11 downto 2);
					when 304 => temp(3049 downto 3040) := ADC(11 downto 2);
					when 305 => temp(3059 downto 3050) := ADC(11 downto 2);
					when 306 => temp(3069 downto 3060) := ADC(11 downto 2);
					when 307 => temp(3079 downto 3070) := ADC(11 downto 2);
					when 308 => temp(3089 downto 3080) := ADC(11 downto 2);
					when 309 => temp(3099 downto 3090) := ADC(11 downto 2);
					when 310 => temp(3109 downto 3100) := ADC(11 downto 2);
					when 311 => temp(3119 downto 3110) := ADC(11 downto 2);
					when 312 => temp(3129 downto 3120) := ADC(11 downto 2);
					when 313 => temp(3139 downto 3130) := ADC(11 downto 2);
					when 314 => temp(3149 downto 3140) := ADC(11 downto 2);
					when 315 => temp(3159 downto 3150) := ADC(11 downto 2);
					when 316 => temp(3169 downto 3160) := ADC(11 downto 2);
					when 317 => temp(3179 downto 3170) := ADC(11 downto 2);
					when 318 => temp(3189 downto 3180) := ADC(11 downto 2);
					when 319 => temp(3199 downto 3190) := ADC(11 downto 2);
					when 320 => temp(3209 downto 3200) := ADC(11 downto 2);
					when 321 => temp(3219 downto 3210) := ADC(11 downto 2);
					when 322 => temp(3229 downto 3220) := ADC(11 downto 2);
					when 323 => temp(3239 downto 3230) := ADC(11 downto 2);
					when 324 => temp(3249 downto 3240) := ADC(11 downto 2);
					when 325 => temp(3259 downto 3250) := ADC(11 downto 2);
					when 326 => temp(3269 downto 3260) := ADC(11 downto 2);
					when 327 => temp(3279 downto 3270) := ADC(11 downto 2);
					when 328 => temp(3289 downto 3280) := ADC(11 downto 2);
					when 329 => temp(3299 downto 3290) := ADC(11 downto 2);
					when 330 => temp(3309 downto 3300) := ADC(11 downto 2);
					when 331 => temp(3319 downto 3310) := ADC(11 downto 2);
					when 332 => temp(3329 downto 3320) := ADC(11 downto 2);
					when 333 => temp(3339 downto 3330) := ADC(11 downto 2);
					when 334 => temp(3349 downto 3340) := ADC(11 downto 2);
					when 335 => temp(3359 downto 3350) := ADC(11 downto 2);
					when 336 => temp(3369 downto 3360) := ADC(11 downto 2);
					when 337 => temp(3379 downto 3370) := ADC(11 downto 2);
					when 338 => temp(3389 downto 3380) := ADC(11 downto 2);
					when 339 => temp(3399 downto 3390) := ADC(11 downto 2);
					when 340 => temp(3409 downto 3400) := ADC(11 downto 2);
					when 341 => temp(3419 downto 3410) := ADC(11 downto 2);
					when 342 => temp(3429 downto 3420) := ADC(11 downto 2);
					when 343 => temp(3439 downto 3430) := ADC(11 downto 2);
					when 344 => temp(3449 downto 3440) := ADC(11 downto 2);
					when 345 => temp(3459 downto 3450) := ADC(11 downto 2);
					when 346 => temp(3469 downto 3460) := ADC(11 downto 2);
					when 347 => temp(3479 downto 3470) := ADC(11 downto 2);
					when 348 => temp(3489 downto 3480) := ADC(11 downto 2);
					when 349 => temp(3499 downto 3490) := ADC(11 downto 2);
					when 350 => temp(3509 downto 3500) := ADC(11 downto 2);
					when 351 => temp(3519 downto 3510) := ADC(11 downto 2);
					when 352 => temp(3529 downto 3520) := ADC(11 downto 2);
					when 353 => temp(3539 downto 3530) := ADC(11 downto 2);
					when 354 => temp(3549 downto 3540) := ADC(11 downto 2);
					when 355 => temp(3559 downto 3550) := ADC(11 downto 2);
					when 356 => temp(3569 downto 3560) := ADC(11 downto 2);
					when 357 => temp(3579 downto 3570) := ADC(11 downto 2);
					when 358 => temp(3589 downto 3580) := ADC(11 downto 2);
					when 359 => temp(3599 downto 3590) := ADC(11 downto 2);
					when 360 => temp(3609 downto 3600) := ADC(11 downto 2);
					when 361 => temp(3619 downto 3610) := ADC(11 downto 2);
					when 362 => temp(3629 downto 3620) := ADC(11 downto 2);
					when 363 => temp(3639 downto 3630) := ADC(11 downto 2);
					when 364 => temp(3649 downto 3640) := ADC(11 downto 2);
					when 365 => temp(3659 downto 3650) := ADC(11 downto 2);
					when 366 => temp(3669 downto 3660) := ADC(11 downto 2);
					when 367 => temp(3679 downto 3670) := ADC(11 downto 2);
					when 368 => temp(3689 downto 3680) := ADC(11 downto 2);
					when 369 => temp(3699 downto 3690) := ADC(11 downto 2);
					when 370 => temp(3709 downto 3700) := ADC(11 downto 2);
					when 371 => temp(3719 downto 3710) := ADC(11 downto 2);
					when 372 => temp(3729 downto 3720) := ADC(11 downto 2);
					when 373 => temp(3739 downto 3730) := ADC(11 downto 2);
					when 374 => temp(3749 downto 3740) := ADC(11 downto 2);
					when 375 => temp(3759 downto 3750) := ADC(11 downto 2);
					when 376 => temp(3769 downto 3760) := ADC(11 downto 2);
					when 377 => temp(3779 downto 3770) := ADC(11 downto 2);
					when 378 => temp(3789 downto 3780) := ADC(11 downto 2);
					when 379 => temp(3799 downto 3790) := ADC(11 downto 2);
					when 380 => temp(3809 downto 3800) := ADC(11 downto 2);
					when 381 => temp(3819 downto 3810) := ADC(11 downto 2);
					when 382 => temp(3829 downto 3820) := ADC(11 downto 2);
					when 383 => temp(3839 downto 3830) := ADC(11 downto 2);
					when 384 => temp(3849 downto 3840) := ADC(11 downto 2);
					when 385 => temp(3859 downto 3850) := ADC(11 downto 2);
					when 386 => temp(3869 downto 3860) := ADC(11 downto 2);
					when 387 => temp(3879 downto 3870) := ADC(11 downto 2);
					when 388 => temp(3889 downto 3880) := ADC(11 downto 2);
					when 389 => temp(3899 downto 3890) := ADC(11 downto 2);
					when 390 => temp(3909 downto 3900) := ADC(11 downto 2);
					when 391 => temp(3919 downto 3910) := ADC(11 downto 2);
					when 392 => temp(3929 downto 3920) := ADC(11 downto 2);
					when 393 => temp(3939 downto 3930) := ADC(11 downto 2);
					when 394 => temp(3949 downto 3940) := ADC(11 downto 2);
					when 395 => temp(3959 downto 3950) := ADC(11 downto 2);
					when 396 => temp(3969 downto 3960) := ADC(11 downto 2);
					when 397 => temp(3979 downto 3970) := ADC(11 downto 2);
					when 398 => temp(3989 downto 3980) := ADC(11 downto 2);
					when 399 => temp(3999 downto 3990) := ADC(11 downto 2);
					when 400 => temp(4009 downto 4000) := ADC(11 downto 2);
					when 401 => temp(4019 downto 4010) := ADC(11 downto 2);
					when 402 => temp(4029 downto 4020) := ADC(11 downto 2);
					when 403 => temp(4039 downto 4030) := ADC(11 downto 2);
					when 404 => temp(4049 downto 4040) := ADC(11 downto 2);
					when 405 => temp(4059 downto 4050) := ADC(11 downto 2);
					when 406 => temp(4069 downto 4060) := ADC(11 downto 2);
					when 407 => temp(4079 downto 4070) := ADC(11 downto 2);
					when 408 => temp(4089 downto 4080) := ADC(11 downto 2);
					when 409 => temp(4099 downto 4090) := ADC(11 downto 2);
					when 410 => temp(4109 downto 4100) := ADC(11 downto 2);
					when 411 => temp(4119 downto 4110) := ADC(11 downto 2);
					when 412 => temp(4129 downto 4120) := ADC(11 downto 2);
					when 413 => temp(4139 downto 4130) := ADC(11 downto 2);
					when 414 => temp(4149 downto 4140) := ADC(11 downto 2);
					when 415 => temp(4159 downto 4150) := ADC(11 downto 2);
					when 416 => temp(4169 downto 4160) := ADC(11 downto 2);
					when 417 => temp(4179 downto 4170) := ADC(11 downto 2);
					when 418 => temp(4189 downto 4180) := ADC(11 downto 2);
					when 419 => temp(4199 downto 4190) := ADC(11 downto 2);
					when 420 => temp(4209 downto 4200) := ADC(11 downto 2);
					when 421 => temp(4219 downto 4210) := ADC(11 downto 2);
					when 422 => temp(4229 downto 4220) := ADC(11 downto 2);
					when 423 => temp(4239 downto 4230) := ADC(11 downto 2);
					when 424 => temp(4249 downto 4240) := ADC(11 downto 2);
					when 425 => temp(4259 downto 4250) := ADC(11 downto 2);
					when 426 => temp(4269 downto 4260) := ADC(11 downto 2);
					when 427 => temp(4279 downto 4270) := ADC(11 downto 2);
					when 428 => temp(4289 downto 4280) := ADC(11 downto 2);
					when 429 => temp(4299 downto 4290) := ADC(11 downto 2);
					when 430 => temp(4309 downto 4300) := ADC(11 downto 2);
					when 431 => temp(4319 downto 4310) := ADC(11 downto 2);
					when 432 => temp(4329 downto 4320) := ADC(11 downto 2);
					when 433 => temp(4339 downto 4330) := ADC(11 downto 2);
					when 434 => temp(4349 downto 4340) := ADC(11 downto 2);
					when 435 => temp(4359 downto 4350) := ADC(11 downto 2);
					when 436 => temp(4369 downto 4360) := ADC(11 downto 2);
					when 437 => temp(4379 downto 4370) := ADC(11 downto 2);
					when 438 => temp(4389 downto 4380) := ADC(11 downto 2);
					when 439 => temp(4399 downto 4390) := ADC(11 downto 2);
					when 440 => temp(4409 downto 4400) := ADC(11 downto 2);
					when 441 => temp(4419 downto 4410) := ADC(11 downto 2);
					when 442 => temp(4429 downto 4420) := ADC(11 downto 2);
					when 443 => temp(4439 downto 4430) := ADC(11 downto 2);
					when 444 => temp(4449 downto 4440) := ADC(11 downto 2);
					when 445 => temp(4459 downto 4450) := ADC(11 downto 2);
					when 446 => temp(4469 downto 4460) := ADC(11 downto 2);
					when 447 => temp(4479 downto 4470) := ADC(11 downto 2);
					when 448 => temp(4489 downto 4480) := ADC(11 downto 2);
					when 449 => temp(4499 downto 4490) := ADC(11 downto 2);
					when 450 => temp(4509 downto 4500) := ADC(11 downto 2);
					when 451 => temp(4519 downto 4510) := ADC(11 downto 2);
					when 452 => temp(4529 downto 4520) := ADC(11 downto 2);
					when 453 => temp(4539 downto 4530) := ADC(11 downto 2);
					when 454 => temp(4549 downto 4540) := ADC(11 downto 2);
					when 455 => temp(4559 downto 4550) := ADC(11 downto 2);
					when 456 => temp(4569 downto 4560) := ADC(11 downto 2);
					when 457 => temp(4579 downto 4570) := ADC(11 downto 2);
					when 458 => temp(4589 downto 4580) := ADC(11 downto 2);
					when 459 => temp(4599 downto 4590) := ADC(11 downto 2);
					when 460 => temp(4609 downto 4600) := ADC(11 downto 2);
					when 461 => temp(4619 downto 4610) := ADC(11 downto 2);
					when 462 => temp(4629 downto 4620) := ADC(11 downto 2);
					when 463 => temp(4639 downto 4630) := ADC(11 downto 2);
					when 464 => temp(4649 downto 4640) := ADC(11 downto 2);
					when 465 => temp(4659 downto 4650) := ADC(11 downto 2);
					when 466 => temp(4669 downto 4660) := ADC(11 downto 2);
					when 467 => temp(4679 downto 4670) := ADC(11 downto 2);
					when 468 => temp(4689 downto 4680) := ADC(11 downto 2);
					when 469 => temp(4699 downto 4690) := ADC(11 downto 2);
					when 470 => temp(4709 downto 4700) := ADC(11 downto 2);
					when 471 => temp(4719 downto 4710) := ADC(11 downto 2);
					when 472 => temp(4729 downto 4720) := ADC(11 downto 2);
					when 473 => temp(4739 downto 4730) := ADC(11 downto 2);
					when 474 => temp(4749 downto 4740) := ADC(11 downto 2);
					when 475 => temp(4759 downto 4750) := ADC(11 downto 2);
					when 476 => temp(4769 downto 4760) := ADC(11 downto 2);
					when 477 => temp(4779 downto 4770) := ADC(11 downto 2);
					when 478 => temp(4789 downto 4780) := ADC(11 downto 2);
					when 479 => temp(4799 downto 4790) := ADC(11 downto 2);
					when 480 => temp(4809 downto 4800) := ADC(11 downto 2);
					when 481 => temp(4819 downto 4810) := ADC(11 downto 2);
					when 482 => temp(4829 downto 4820) := ADC(11 downto 2);
					when 483 => temp(4839 downto 4830) := ADC(11 downto 2);
					when 484 => temp(4849 downto 4840) := ADC(11 downto 2);
					when 485 => temp(4859 downto 4850) := ADC(11 downto 2);
					when 486 => temp(4869 downto 4860) := ADC(11 downto 2);
					when 487 => temp(4879 downto 4870) := ADC(11 downto 2);
					when 488 => temp(4889 downto 4880) := ADC(11 downto 2);
					when 489 => temp(4899 downto 4890) := ADC(11 downto 2);
					when 490 => temp(4909 downto 4900) := ADC(11 downto 2);
					when 491 => temp(4919 downto 4910) := ADC(11 downto 2);
					when 492 => temp(4929 downto 4920) := ADC(11 downto 2);
					when 493 => temp(4939 downto 4930) := ADC(11 downto 2);
					when 494 => temp(4949 downto 4940) := ADC(11 downto 2);
					when 495 => temp(4959 downto 4950) := ADC(11 downto 2);
					when 496 => temp(4969 downto 4960) := ADC(11 downto 2);
					when 497 => temp(4979 downto 4970) := ADC(11 downto 2);
					when 498 => temp(4989 downto 4980) := ADC(11 downto 2);
					when 499 => temp(4999 downto 4990) := ADC(11 downto 2);
					when 500 => temp(5009 downto 5000) := ADC(11 downto 2);
					when 501 => temp(5019 downto 5010) := ADC(11 downto 2);
					when 502 => temp(5029 downto 5020) := ADC(11 downto 2);
					when 503 => temp(5039 downto 5030) := ADC(11 downto 2);
					when 504 => temp(5049 downto 5040) := ADC(11 downto 2);
					when 505 => temp(5059 downto 5050) := ADC(11 downto 2);
					when 506 => temp(5069 downto 5060) := ADC(11 downto 2);
					when 507 => temp(5079 downto 5070) := ADC(11 downto 2);
					when 508 => temp(5089 downto 5080) := ADC(11 downto 2);
					when 509 => temp(5099 downto 5090) := ADC(11 downto 2);
					when 510 => temp(5109 downto 5100) := ADC(11 downto 2);
					when 511 => temp(5119 downto 5110) := ADC(11 downto 2);
					when 512 => temp(5129 downto 5120) := ADC(11 downto 2);
					when 513 => temp(5139 downto 5130) := ADC(11 downto 2);
					when 514 => temp(5149 downto 5140) := ADC(11 downto 2);
					when 515 => temp(5159 downto 5150) := ADC(11 downto 2);
					when 516 => temp(5169 downto 5160) := ADC(11 downto 2);
					when 517 => temp(5179 downto 5170) := ADC(11 downto 2);
					when 518 => temp(5189 downto 5180) := ADC(11 downto 2);
					when 519 => temp(5199 downto 5190) := ADC(11 downto 2);
					when 520 => temp(5209 downto 5200) := ADC(11 downto 2);
					when 521 => temp(5219 downto 5210) := ADC(11 downto 2);
					when 522 => temp(5229 downto 5220) := ADC(11 downto 2);
					when 523 => temp(5239 downto 5230) := ADC(11 downto 2);
					when 524 => temp(5249 downto 5240) := ADC(11 downto 2);
					when 525 => temp(5259 downto 5250) := ADC(11 downto 2);
					when 526 => temp(5269 downto 5260) := ADC(11 downto 2);
					when 527 => temp(5279 downto 5270) := ADC(11 downto 2);
					when 528 => temp(5289 downto 5280) := ADC(11 downto 2);
					when 529 => temp(5299 downto 5290) := ADC(11 downto 2);
					when 530 => temp(5309 downto 5300) := ADC(11 downto 2);
					when 531 => temp(5319 downto 5310) := ADC(11 downto 2);
					when 532 => temp(5329 downto 5320) := ADC(11 downto 2);
					when 533 => temp(5339 downto 5330) := ADC(11 downto 2);
					when 534 => temp(5349 downto 5340) := ADC(11 downto 2);
					when 535 => temp(5359 downto 5350) := ADC(11 downto 2);
					when 536 => temp(5369 downto 5360) := ADC(11 downto 2);
					when 537 => temp(5379 downto 5370) := ADC(11 downto 2);
					when 538 => temp(5389 downto 5380) := ADC(11 downto 2);
					when 539 => temp(5399 downto 5390) := ADC(11 downto 2);
					when 540 => temp(5409 downto 5400) := ADC(11 downto 2);
					when 541 => temp(5419 downto 5410) := ADC(11 downto 2);
					when 542 => temp(5429 downto 5420) := ADC(11 downto 2);
					when 543 => temp(5439 downto 5430) := ADC(11 downto 2);
					when 544 => temp(5449 downto 5440) := ADC(11 downto 2);
					when 545 => temp(5459 downto 5450) := ADC(11 downto 2);
					when 546 => temp(5469 downto 5460) := ADC(11 downto 2);
					when 547 => temp(5479 downto 5470) := ADC(11 downto 2);
					when 548 => temp(5489 downto 5480) := ADC(11 downto 2);
					when 549 => temp(5499 downto 5490) := ADC(11 downto 2);
					when 550 => temp(5509 downto 5500) := ADC(11 downto 2);
					when 551 => temp(5519 downto 5510) := ADC(11 downto 2);
					when 552 => temp(5529 downto 5520) := ADC(11 downto 2);
					when 553 => temp(5539 downto 5530) := ADC(11 downto 2);
					when 554 => temp(5549 downto 5540) := ADC(11 downto 2);
					when 555 => temp(5559 downto 5550) := ADC(11 downto 2);
					when 556 => temp(5569 downto 5560) := ADC(11 downto 2);
					when 557 => temp(5579 downto 5570) := ADC(11 downto 2);
					when 558 => temp(5589 downto 5580) := ADC(11 downto 2);
					when 559 => temp(5599 downto 5590) := ADC(11 downto 2);
					when 560 => temp(5609 downto 5600) := ADC(11 downto 2);
					when 561 => temp(5619 downto 5610) := ADC(11 downto 2);
					when 562 => temp(5629 downto 5620) := ADC(11 downto 2);
					when 563 => temp(5639 downto 5630) := ADC(11 downto 2);
					when 564 => temp(5649 downto 5640) := ADC(11 downto 2);
					when 565 => temp(5659 downto 5650) := ADC(11 downto 2);
					when 566 => temp(5669 downto 5660) := ADC(11 downto 2);
					when 567 => temp(5679 downto 5670) := ADC(11 downto 2);
					when 568 => temp(5689 downto 5680) := ADC(11 downto 2);
					when 569 => temp(5699 downto 5690) := ADC(11 downto 2);
					when 570 => temp(5709 downto 5700) := ADC(11 downto 2);
					when 571 => temp(5719 downto 5710) := ADC(11 downto 2);
					when 572 => temp(5729 downto 5720) := ADC(11 downto 2);
					when 573 => temp(5739 downto 5730) := ADC(11 downto 2);
					when 574 => temp(5749 downto 5740) := ADC(11 downto 2);
					when 575 => temp(5759 downto 5750) := ADC(11 downto 2);
					when 576 => temp(5769 downto 5760) := ADC(11 downto 2);
					when 577 => temp(5779 downto 5770) := ADC(11 downto 2);
					when 578 => temp(5789 downto 5780) := ADC(11 downto 2);
					when 579 => temp(5799 downto 5790) := ADC(11 downto 2);
					when 580 => temp(5809 downto 5800) := ADC(11 downto 2);
					when 581 => temp(5819 downto 5810) := ADC(11 downto 2);
					when 582 => temp(5829 downto 5820) := ADC(11 downto 2);
					when 583 => temp(5839 downto 5830) := ADC(11 downto 2);
					when 584 => temp(5849 downto 5840) := ADC(11 downto 2);
					when 585 => temp(5859 downto 5850) := ADC(11 downto 2);
					when 586 => temp(5869 downto 5860) := ADC(11 downto 2);
					when 587 => temp(5879 downto 5870) := ADC(11 downto 2);
					when 588 => temp(5889 downto 5880) := ADC(11 downto 2);
					when 589 => temp(5899 downto 5890) := ADC(11 downto 2);
					when 590 => temp(5909 downto 5900) := ADC(11 downto 2);
					when 591 => temp(5919 downto 5910) := ADC(11 downto 2);
					when 592 => temp(5929 downto 5920) := ADC(11 downto 2);
					when 593 => temp(5939 downto 5930) := ADC(11 downto 2);
					when 594 => temp(5949 downto 5940) := ADC(11 downto 2);
					when 595 => temp(5959 downto 5950) := ADC(11 downto 2);
					when 596 => temp(5969 downto 5960) := ADC(11 downto 2);
					when 597 => temp(5979 downto 5970) := ADC(11 downto 2);
					when 598 => temp(5989 downto 5980) := ADC(11 downto 2);
					when 599 => temp(5999 downto 5990) := ADC(11 downto 2);
					when 600 => temp(6009 downto 6000) := ADC(11 downto 2);
					when 601 => temp(6019 downto 6010) := ADC(11 downto 2);
					when 602 => temp(6029 downto 6020) := ADC(11 downto 2);
					when 603 => temp(6039 downto 6030) := ADC(11 downto 2);
					when 604 => temp(6049 downto 6040) := ADC(11 downto 2);
					when 605 => temp(6059 downto 6050) := ADC(11 downto 2);
					when 606 => temp(6069 downto 6060) := ADC(11 downto 2);
					when 607 => temp(6079 downto 6070) := ADC(11 downto 2);
					when 608 => temp(6089 downto 6080) := ADC(11 downto 2);
					when 609 => temp(6099 downto 6090) := ADC(11 downto 2);
					when 610 => temp(6109 downto 6100) := ADC(11 downto 2);
					when 611 => temp(6119 downto 6110) := ADC(11 downto 2);
					when 612 => temp(6129 downto 6120) := ADC(11 downto 2);
					when 613 => temp(6139 downto 6130) := ADC(11 downto 2);
					when 614 => temp(6149 downto 6140) := ADC(11 downto 2);
					when 615 => temp(6159 downto 6150) := ADC(11 downto 2);
					when 616 => temp(6169 downto 6160) := ADC(11 downto 2);
					when 617 => temp(6179 downto 6170) := ADC(11 downto 2);
					when 618 => temp(6189 downto 6180) := ADC(11 downto 2);
					when 619 => temp(6199 downto 6190) := ADC(11 downto 2);
					when 620 => temp(6209 downto 6200) := ADC(11 downto 2);
					when 621 => temp(6219 downto 6210) := ADC(11 downto 2);
					when 622 => temp(6229 downto 6220) := ADC(11 downto 2);
					when 623 => temp(6239 downto 6230) := ADC(11 downto 2);
					when 624 => temp(6249 downto 6240) := ADC(11 downto 2);
					when 625 => temp(6259 downto 6250) := ADC(11 downto 2);
					when 626 => temp(6269 downto 6260) := ADC(11 downto 2);
					when 627 => temp(6279 downto 6270) := ADC(11 downto 2);
					when 628 => temp(6289 downto 6280) := ADC(11 downto 2);
					when 629 => temp(6299 downto 6290) := ADC(11 downto 2);
					when 630 => temp(6309 downto 6300) := ADC(11 downto 2);
					when 631 => temp(6319 downto 6310) := ADC(11 downto 2);
					when 632 => temp(6329 downto 6320) := ADC(11 downto 2);
					when 633 => temp(6339 downto 6330) := ADC(11 downto 2);
					when 634 => temp(6349 downto 6340) := ADC(11 downto 2);
					when 635 => temp(6359 downto 6350) := ADC(11 downto 2);
					when 636 => temp(6369 downto 6360) := ADC(11 downto 2);
					when 637 => temp(6379 downto 6370) := ADC(11 downto 2);
					when 638 => temp(6389 downto 6380) := ADC(11 downto 2);
					when 639 => temp(6399 downto 6390) := ADC(11 downto 2);
					when 640 => temp(6409 downto 6400) := ADC(11 downto 2);
					when 641 => temp(6419 downto 6410) := ADC(11 downto 2);
					when 642 => temp(6429 downto 6420) := ADC(11 downto 2);
					when 643 => temp(6439 downto 6430) := ADC(11 downto 2);
					when 644 => temp(6449 downto 6440) := ADC(11 downto 2);
					when 645 => temp(6459 downto 6450) := ADC(11 downto 2);
					when 646 => temp(6469 downto 6460) := ADC(11 downto 2);
					when 647 => temp(6479 downto 6470) := ADC(11 downto 2);
					when 648 => temp(6489 downto 6480) := ADC(11 downto 2);
					when 649 => temp(6499 downto 6490) := ADC(11 downto 2);
					when 650 => temp(6509 downto 6500) := ADC(11 downto 2);
					when 651 => temp(6519 downto 6510) := ADC(11 downto 2);
					when 652 => temp(6529 downto 6520) := ADC(11 downto 2);
					when 653 => temp(6539 downto 6530) := ADC(11 downto 2);
					when 654 => temp(6549 downto 6540) := ADC(11 downto 2);
					when 655 => temp(6559 downto 6550) := ADC(11 downto 2);
					when 656 => temp(6569 downto 6560) := ADC(11 downto 2);
					when 657 => temp(6579 downto 6570) := ADC(11 downto 2);
					when 658 => temp(6589 downto 6580) := ADC(11 downto 2);
					when 659 => temp(6599 downto 6590) := ADC(11 downto 2);
					when 660 => temp(6609 downto 6600) := ADC(11 downto 2);
					when 661 => temp(6619 downto 6610) := ADC(11 downto 2);
					when 662 => temp(6629 downto 6620) := ADC(11 downto 2);
					when 663 => temp(6639 downto 6630) := ADC(11 downto 2);
					when 664 => temp(6649 downto 6640) := ADC(11 downto 2);
					when 665 => temp(6659 downto 6650) := ADC(11 downto 2);
					when 666 => temp(6669 downto 6660) := ADC(11 downto 2);
					when 667 => temp(6679 downto 6670) := ADC(11 downto 2);
					when 668 => temp(6689 downto 6680) := ADC(11 downto 2);
					when 669 => temp(6699 downto 6690) := ADC(11 downto 2);
					when 670 => temp(6709 downto 6700) := ADC(11 downto 2);
					when 671 => temp(6719 downto 6710) := ADC(11 downto 2);
					when 672 => temp(6729 downto 6720) := ADC(11 downto 2);
					when 673 => temp(6739 downto 6730) := ADC(11 downto 2);
					when 674 => temp(6749 downto 6740) := ADC(11 downto 2);
					when 675 => temp(6759 downto 6750) := ADC(11 downto 2);
					when 676 => temp(6769 downto 6760) := ADC(11 downto 2);
					when 677 => temp(6779 downto 6770) := ADC(11 downto 2);
					when 678 => temp(6789 downto 6780) := ADC(11 downto 2);
					when 679 => temp(6799 downto 6790) := ADC(11 downto 2);
					when 680 => temp(6809 downto 6800) := ADC(11 downto 2);
					when 681 => temp(6819 downto 6810) := ADC(11 downto 2);
					when 682 => temp(6829 downto 6820) := ADC(11 downto 2);
					when 683 => temp(6839 downto 6830) := ADC(11 downto 2);
					when 684 => temp(6849 downto 6840) := ADC(11 downto 2);
					when 685 => temp(6859 downto 6850) := ADC(11 downto 2);
					when 686 => temp(6869 downto 6860) := ADC(11 downto 2);
					when 687 => temp(6879 downto 6870) := ADC(11 downto 2);
					when 688 => temp(6889 downto 6880) := ADC(11 downto 2);
					when 689 => temp(6899 downto 6890) := ADC(11 downto 2);
					when 690 => temp(6909 downto 6900) := ADC(11 downto 2);
					when 691 => temp(6919 downto 6910) := ADC(11 downto 2);
					when 692 => temp(6929 downto 6920) := ADC(11 downto 2);
					when 693 => temp(6939 downto 6930) := ADC(11 downto 2);
					when 694 => temp(6949 downto 6940) := ADC(11 downto 2);
					when 695 => temp(6959 downto 6950) := ADC(11 downto 2);
					when 696 => temp(6969 downto 6960) := ADC(11 downto 2);
					when 697 => temp(6979 downto 6970) := ADC(11 downto 2);
					when 698 => temp(6989 downto 6980) := ADC(11 downto 2);
					when 699 => temp(6999 downto 6990) := ADC(11 downto 2);
					when 700 => temp(7009 downto 7000) := ADC(11 downto 2);
					when 701 => temp(7019 downto 7010) := ADC(11 downto 2);
					when 702 => temp(7029 downto 7020) := ADC(11 downto 2);
					when 703 => temp(7039 downto 7030) := ADC(11 downto 2);
					when 704 => temp(7049 downto 7040) := ADC(11 downto 2);
					when 705 => temp(7059 downto 7050) := ADC(11 downto 2);
					when 706 => temp(7069 downto 7060) := ADC(11 downto 2);
					when 707 => temp(7079 downto 7070) := ADC(11 downto 2);
					when 708 => temp(7089 downto 7080) := ADC(11 downto 2);
					when 709 => temp(7099 downto 7090) := ADC(11 downto 2);
					when 710 => temp(7109 downto 7100) := ADC(11 downto 2);
					when 711 => temp(7119 downto 7110) := ADC(11 downto 2);
					when 712 => temp(7129 downto 7120) := ADC(11 downto 2);
					when 713 => temp(7139 downto 7130) := ADC(11 downto 2);
					when 714 => temp(7149 downto 7140) := ADC(11 downto 2);
					when 715 => temp(7159 downto 7150) := ADC(11 downto 2);
					when 716 => temp(7169 downto 7160) := ADC(11 downto 2);
					when 717 => temp(7179 downto 7170) := ADC(11 downto 2);
					when 718 => temp(7189 downto 7180) := ADC(11 downto 2);
					when 719 => temp(7199 downto 7190) := ADC(11 downto 2);
					when 720 => temp(7209 downto 7200) := ADC(11 downto 2);
					when 721 => temp(7219 downto 7210) := ADC(11 downto 2);
					when 722 => temp(7229 downto 7220) := ADC(11 downto 2);
					when 723 => temp(7239 downto 7230) := ADC(11 downto 2);
					when 724 => temp(7249 downto 7240) := ADC(11 downto 2);
					when 725 => temp(7259 downto 7250) := ADC(11 downto 2);
					when 726 => temp(7269 downto 7260) := ADC(11 downto 2);
					when 727 => temp(7279 downto 7270) := ADC(11 downto 2);
					when 728 => temp(7289 downto 7280) := ADC(11 downto 2);
					when 729 => temp(7299 downto 7290) := ADC(11 downto 2);
					when 730 => temp(7309 downto 7300) := ADC(11 downto 2);
					when 731 => temp(7319 downto 7310) := ADC(11 downto 2);
					when 732 => temp(7329 downto 7320) := ADC(11 downto 2);
					when 733 => temp(7339 downto 7330) := ADC(11 downto 2);
					when 734 => temp(7349 downto 7340) := ADC(11 downto 2);
					when 735 => temp(7359 downto 7350) := ADC(11 downto 2);
					when 736 => temp(7369 downto 7360) := ADC(11 downto 2);
					when 737 => temp(7379 downto 7370) := ADC(11 downto 2);
					when 738 => temp(7389 downto 7380) := ADC(11 downto 2);
					when 739 => temp(7399 downto 7390) := ADC(11 downto 2);
					when 740 => temp(7409 downto 7400) := ADC(11 downto 2);
					when 741 => temp(7419 downto 7410) := ADC(11 downto 2);
					when 742 => temp(7429 downto 7420) := ADC(11 downto 2);
					when 743 => temp(7439 downto 7430) := ADC(11 downto 2);
					when 744 => temp(7449 downto 7440) := ADC(11 downto 2);
					when 745 => temp(7459 downto 7450) := ADC(11 downto 2);
					when 746 => temp(7469 downto 7460) := ADC(11 downto 2);
					when 747 => temp(7479 downto 7470) := ADC(11 downto 2);
					when 748 => temp(7489 downto 7480) := ADC(11 downto 2);
					when 749 => temp(7499 downto 7490) := ADC(11 downto 2);
					when 750 => temp(7509 downto 7500) := ADC(11 downto 2);
					when 751 => temp(7519 downto 7510) := ADC(11 downto 2);
					when 752 => temp(7529 downto 7520) := ADC(11 downto 2);
					when 753 => temp(7539 downto 7530) := ADC(11 downto 2);
					when 754 => temp(7549 downto 7540) := ADC(11 downto 2);
					when 755 => temp(7559 downto 7550) := ADC(11 downto 2);
					when 756 => temp(7569 downto 7560) := ADC(11 downto 2);
					when 757 => temp(7579 downto 7570) := ADC(11 downto 2);
					when 758 => temp(7589 downto 7580) := ADC(11 downto 2);
					when 759 => temp(7599 downto 7590) := ADC(11 downto 2);
					when 760 => temp(7609 downto 7600) := ADC(11 downto 2);
					when 761 => temp(7619 downto 7610) := ADC(11 downto 2);
					when 762 => temp(7629 downto 7620) := ADC(11 downto 2);
					when 763 => temp(7639 downto 7630) := ADC(11 downto 2);
					when 764 => temp(7649 downto 7640) := ADC(11 downto 2);
					when 765 => temp(7659 downto 7650) := ADC(11 downto 2);
					when 766 => temp(7669 downto 7660) := ADC(11 downto 2);
					when 767 => temp(7679 downto 7670) := ADC(11 downto 2);
					when 768 => temp(7689 downto 7680) := ADC(11 downto 2);
					when 769 => temp(7699 downto 7690) := ADC(11 downto 2);
					when 770 => temp(7709 downto 7700) := ADC(11 downto 2);
					when 771 => temp(7719 downto 7710) := ADC(11 downto 2);
					when 772 => temp(7729 downto 7720) := ADC(11 downto 2);
					when 773 => temp(7739 downto 7730) := ADC(11 downto 2);
					when 774 => temp(7749 downto 7740) := ADC(11 downto 2);
					when 775 => temp(7759 downto 7750) := ADC(11 downto 2);
					when 776 => temp(7769 downto 7760) := ADC(11 downto 2);
					when 777 => temp(7779 downto 7770) := ADC(11 downto 2);
					when 778 => temp(7789 downto 7780) := ADC(11 downto 2);
					when 779 => temp(7799 downto 7790) := ADC(11 downto 2);
					when 780 => temp(7809 downto 7800) := ADC(11 downto 2);
					when 781 => temp(7819 downto 7810) := ADC(11 downto 2);
					when 782 => temp(7829 downto 7820) := ADC(11 downto 2);
					when 783 => temp(7839 downto 7830) := ADC(11 downto 2);
					when 784 => temp(7849 downto 7840) := ADC(11 downto 2);
					when 785 => temp(7859 downto 7850) := ADC(11 downto 2);
					when 786 => temp(7869 downto 7860) := ADC(11 downto 2);
					when 787 => temp(7879 downto 7870) := ADC(11 downto 2);
					when 788 => temp(7889 downto 7880) := ADC(11 downto 2);
					when 789 => temp(7899 downto 7890) := ADC(11 downto 2);
					when 790 => temp(7909 downto 7900) := ADC(11 downto 2);
					when 791 => temp(7919 downto 7910) := ADC(11 downto 2);
					when 792 => temp(7929 downto 7920) := ADC(11 downto 2);
					when 793 => temp(7939 downto 7930) := ADC(11 downto 2);
					when 794 => temp(7949 downto 7940) := ADC(11 downto 2);
					when 795 => temp(7959 downto 7950) := ADC(11 downto 2);
					when 796 => temp(7969 downto 7960) := ADC(11 downto 2);
					when 797 => temp(7979 downto 7970) := ADC(11 downto 2);
					when 798 => temp(7989 downto 7980) := ADC(11 downto 2);
					when 799 => temp(7999 downto 7990) := ADC(11 downto 2);
					when 800 => temp(8009 downto 8000) := ADC(11 downto 2);
					when 801 => temp(8019 downto 8010) := ADC(11 downto 2);
					when 802 => temp(8029 downto 8020) := ADC(11 downto 2);
					when 803 => temp(8039 downto 8030) := ADC(11 downto 2);
					when 804 => temp(8049 downto 8040) := ADC(11 downto 2);
					when 805 => temp(8059 downto 8050) := ADC(11 downto 2);
					when 806 => temp(8069 downto 8060) := ADC(11 downto 2);
					when 807 => temp(8079 downto 8070) := ADC(11 downto 2);
					when 808 => temp(8089 downto 8080) := ADC(11 downto 2);
					when 809 => temp(8099 downto 8090) := ADC(11 downto 2);
					when 810 => temp(8109 downto 8100) := ADC(11 downto 2);
					when 811 => temp(8119 downto 8110) := ADC(11 downto 2);
					when 812 => temp(8129 downto 8120) := ADC(11 downto 2);
					when 813 => temp(8139 downto 8130) := ADC(11 downto 2);
					when 814 => temp(8149 downto 8140) := ADC(11 downto 2);
					when 815 => temp(8159 downto 8150) := ADC(11 downto 2);
					when 816 => temp(8169 downto 8160) := ADC(11 downto 2);
					when 817 => temp(8179 downto 8170) := ADC(11 downto 2);
					when 818 => temp(8189 downto 8180) := ADC(11 downto 2);
					when 819 => temp(8199 downto 8190) := ADC(11 downto 2);
					when 820 => temp(8209 downto 8200) := ADC(11 downto 2);
					when 821 => temp(8219 downto 8210) := ADC(11 downto 2);
					when 822 => temp(8229 downto 8220) := ADC(11 downto 2);
					when 823 => temp(8239 downto 8230) := ADC(11 downto 2);
					when 824 => temp(8249 downto 8240) := ADC(11 downto 2);
					when 825 => temp(8259 downto 8250) := ADC(11 downto 2);
					when 826 => temp(8269 downto 8260) := ADC(11 downto 2);
					when 827 => temp(8279 downto 8270) := ADC(11 downto 2);
					when 828 => temp(8289 downto 8280) := ADC(11 downto 2);
					when 829 => temp(8299 downto 8290) := ADC(11 downto 2);
					when 830 => temp(8309 downto 8300) := ADC(11 downto 2);
					when 831 => temp(8319 downto 8310) := ADC(11 downto 2);
					when 832 => temp(8329 downto 8320) := ADC(11 downto 2);
					when 833 => temp(8339 downto 8330) := ADC(11 downto 2);
					when 834 => temp(8349 downto 8340) := ADC(11 downto 2);
					when 835 => temp(8359 downto 8350) := ADC(11 downto 2);
					when 836 => temp(8369 downto 8360) := ADC(11 downto 2);
					when 837 => temp(8379 downto 8370) := ADC(11 downto 2);
					when 838 => temp(8389 downto 8380) := ADC(11 downto 2);
					when 839 => temp(8399 downto 8390) := ADC(11 downto 2);
					when 840 => temp(8409 downto 8400) := ADC(11 downto 2);
					when 841 => temp(8419 downto 8410) := ADC(11 downto 2);
					when 842 => temp(8429 downto 8420) := ADC(11 downto 2);
					when 843 => temp(8439 downto 8430) := ADC(11 downto 2);
					when 844 => temp(8449 downto 8440) := ADC(11 downto 2);
					when 845 => temp(8459 downto 8450) := ADC(11 downto 2);
					when 846 => temp(8469 downto 8460) := ADC(11 downto 2);
					when 847 => temp(8479 downto 8470) := ADC(11 downto 2);
					when 848 => temp(8489 downto 8480) := ADC(11 downto 2);
					when 849 => temp(8499 downto 8490) := ADC(11 downto 2);
					when 850 => temp(8509 downto 8500) := ADC(11 downto 2);
					when 851 => temp(8519 downto 8510) := ADC(11 downto 2);
					when 852 => temp(8529 downto 8520) := ADC(11 downto 2);
					when 853 => temp(8539 downto 8530) := ADC(11 downto 2);
					when 854 => temp(8549 downto 8540) := ADC(11 downto 2);
					when 855 => temp(8559 downto 8550) := ADC(11 downto 2);
					when 856 => temp(8569 downto 8560) := ADC(11 downto 2);
					when 857 => temp(8579 downto 8570) := ADC(11 downto 2);
					when 858 => temp(8589 downto 8580) := ADC(11 downto 2);
					when 859 => temp(8599 downto 8590) := ADC(11 downto 2);
					when 860 => temp(8609 downto 8600) := ADC(11 downto 2);
					when 861 => temp(8619 downto 8610) := ADC(11 downto 2);
					when 862 => temp(8629 downto 8620) := ADC(11 downto 2);
					when 863 => temp(8639 downto 8630) := ADC(11 downto 2);
					when 864 => temp(8649 downto 8640) := ADC(11 downto 2);
					when 865 => temp(8659 downto 8650) := ADC(11 downto 2);
					when 866 => temp(8669 downto 8660) := ADC(11 downto 2);
					when 867 => temp(8679 downto 8670) := ADC(11 downto 2);
					when 868 => temp(8689 downto 8680) := ADC(11 downto 2);
					when 869 => temp(8699 downto 8690) := ADC(11 downto 2);
					when 870 => temp(8709 downto 8700) := ADC(11 downto 2);
					when 871 => temp(8719 downto 8710) := ADC(11 downto 2);
					when 872 => temp(8729 downto 8720) := ADC(11 downto 2);
					when 873 => temp(8739 downto 8730) := ADC(11 downto 2);
					when 874 => temp(8749 downto 8740) := ADC(11 downto 2);
					when 875 => temp(8759 downto 8750) := ADC(11 downto 2);
					when 876 => temp(8769 downto 8760) := ADC(11 downto 2);
					when 877 => temp(8779 downto 8770) := ADC(11 downto 2);
					when 878 => temp(8789 downto 8780) := ADC(11 downto 2);
					when 879 => temp(8799 downto 8790) := ADC(11 downto 2);
					when 880 => temp(8809 downto 8800) := ADC(11 downto 2);
					when 881 => temp(8819 downto 8810) := ADC(11 downto 2);
					when 882 => temp(8829 downto 8820) := ADC(11 downto 2);
					when 883 => temp(8839 downto 8830) := ADC(11 downto 2);
					when 884 => temp(8849 downto 8840) := ADC(11 downto 2);
					when 885 => temp(8859 downto 8850) := ADC(11 downto 2);
					when 886 => temp(8869 downto 8860) := ADC(11 downto 2);
					when 887 => temp(8879 downto 8870) := ADC(11 downto 2);
					when 888 => temp(8889 downto 8880) := ADC(11 downto 2);
					when 889 => temp(8899 downto 8890) := ADC(11 downto 2);
					when 890 => temp(8909 downto 8900) := ADC(11 downto 2);
					when 891 => temp(8919 downto 8910) := ADC(11 downto 2);
					when 892 => temp(8929 downto 8920) := ADC(11 downto 2);
					when 893 => temp(8939 downto 8930) := ADC(11 downto 2);
					when 894 => temp(8949 downto 8940) := ADC(11 downto 2);
					when 895 => temp(8959 downto 8950) := ADC(11 downto 2);
					when 896 => temp(8969 downto 8960) := ADC(11 downto 2);
					when 897 => temp(8979 downto 8970) := ADC(11 downto 2);
					when 898 => temp(8989 downto 8980) := ADC(11 downto 2);
					when 899 => temp(8999 downto 8990) := ADC(11 downto 2);
					when 900 => temp(9009 downto 9000) := ADC(11 downto 2);
					when 901 => temp(9019 downto 9010) := ADC(11 downto 2);
					when 902 => temp(9029 downto 9020) := ADC(11 downto 2);
					when 903 => temp(9039 downto 9030) := ADC(11 downto 2);
					when 904 => temp(9049 downto 9040) := ADC(11 downto 2);
					when 905 => temp(9059 downto 9050) := ADC(11 downto 2);
					when 906 => temp(9069 downto 9060) := ADC(11 downto 2);
					when 907 => temp(9079 downto 9070) := ADC(11 downto 2);
					when 908 => temp(9089 downto 9080) := ADC(11 downto 2);
					when 909 => temp(9099 downto 9090) := ADC(11 downto 2);
					when 910 => temp(9109 downto 9100) := ADC(11 downto 2);
					when 911 => temp(9119 downto 9110) := ADC(11 downto 2);
					when 912 => temp(9129 downto 9120) := ADC(11 downto 2);
					when 913 => temp(9139 downto 9130) := ADC(11 downto 2);
					when 914 => temp(9149 downto 9140) := ADC(11 downto 2);
					when 915 => temp(9159 downto 9150) := ADC(11 downto 2);
					when 916 => temp(9169 downto 9160) := ADC(11 downto 2);
					when 917 => temp(9179 downto 9170) := ADC(11 downto 2);
					when 918 => temp(9189 downto 9180) := ADC(11 downto 2);
					when 919 => temp(9199 downto 9190) := ADC(11 downto 2);
					when 920 => temp(9209 downto 9200) := ADC(11 downto 2);
					when 921 => temp(9219 downto 9210) := ADC(11 downto 2);
					when 922 => temp(9229 downto 9220) := ADC(11 downto 2);
					when 923 => temp(9239 downto 9230) := ADC(11 downto 2);
					when 924 => temp(9249 downto 9240) := ADC(11 downto 2);
					when 925 => temp(9259 downto 9250) := ADC(11 downto 2);
					when 926 => temp(9269 downto 9260) := ADC(11 downto 2);
					when 927 => temp(9279 downto 9270) := ADC(11 downto 2);
					when 928 => temp(9289 downto 9280) := ADC(11 downto 2);
					when 929 => temp(9299 downto 9290) := ADC(11 downto 2);
					when 930 => temp(9309 downto 9300) := ADC(11 downto 2);
					when 931 => temp(9319 downto 9310) := ADC(11 downto 2);
					when 932 => temp(9329 downto 9320) := ADC(11 downto 2);
					when 933 => temp(9339 downto 9330) := ADC(11 downto 2);
					when 934 => temp(9349 downto 9340) := ADC(11 downto 2);
					when 935 => temp(9359 downto 9350) := ADC(11 downto 2);
					when 936 => temp(9369 downto 9360) := ADC(11 downto 2);
					when 937 => temp(9379 downto 9370) := ADC(11 downto 2);
					when 938 => temp(9389 downto 9380) := ADC(11 downto 2);
					when 939 => temp(9399 downto 9390) := ADC(11 downto 2);
					when 940 => temp(9409 downto 9400) := ADC(11 downto 2);
					when 941 => temp(9419 downto 9410) := ADC(11 downto 2);
					when 942 => temp(9429 downto 9420) := ADC(11 downto 2);
					when 943 => temp(9439 downto 9430) := ADC(11 downto 2);
					when 944 => temp(9449 downto 9440) := ADC(11 downto 2);
					when 945 => temp(9459 downto 9450) := ADC(11 downto 2);
					when 946 => temp(9469 downto 9460) := ADC(11 downto 2);
					when 947 => temp(9479 downto 9470) := ADC(11 downto 2);
					when 948 => temp(9489 downto 9480) := ADC(11 downto 2);
					when 949 => temp(9499 downto 9490) := ADC(11 downto 2);
					when 950 => temp(9509 downto 9500) := ADC(11 downto 2);
					when 951 => temp(9519 downto 9510) := ADC(11 downto 2);
					when 952 => temp(9529 downto 9520) := ADC(11 downto 2);
					when 953 => temp(9539 downto 9530) := ADC(11 downto 2);
					when 954 => temp(9549 downto 9540) := ADC(11 downto 2);
					when 955 => temp(9559 downto 9550) := ADC(11 downto 2);
					when 956 => temp(9569 downto 9560) := ADC(11 downto 2);
					when 957 => temp(9579 downto 9570) := ADC(11 downto 2);
					when 958 => temp(9589 downto 9580) := ADC(11 downto 2);
					when 959 => temp(9599 downto 9590) := ADC(11 downto 2);
					when 960 => temp(9609 downto 9600) := ADC(11 downto 2);
					when 961 => temp(9619 downto 9610) := ADC(11 downto 2);
					when 962 => temp(9629 downto 9620) := ADC(11 downto 2);
					when 963 => temp(9639 downto 9630) := ADC(11 downto 2);
					when 964 => temp(9649 downto 9640) := ADC(11 downto 2);
					when 965 => temp(9659 downto 9650) := ADC(11 downto 2);
					when 966 => temp(9669 downto 9660) := ADC(11 downto 2);
					when 967 => temp(9679 downto 9670) := ADC(11 downto 2);
					when 968 => temp(9689 downto 9680) := ADC(11 downto 2);
					when 969 => temp(9699 downto 9690) := ADC(11 downto 2);
					when 970 => temp(9709 downto 9700) := ADC(11 downto 2);
					when 971 => temp(9719 downto 9710) := ADC(11 downto 2);
					when 972 => temp(9729 downto 9720) := ADC(11 downto 2);
					when 973 => temp(9739 downto 9730) := ADC(11 downto 2);
					when 974 => temp(9749 downto 9740) := ADC(11 downto 2);
					when 975 => temp(9759 downto 9750) := ADC(11 downto 2);
					when 976 => temp(9769 downto 9760) := ADC(11 downto 2);
					when 977 => temp(9779 downto 9770) := ADC(11 downto 2);
					when 978 => temp(9789 downto 9780) := ADC(11 downto 2);
					when 979 => temp(9799 downto 9790) := ADC(11 downto 2);
					when 980 => temp(9809 downto 9800) := ADC(11 downto 2);
					when 981 => temp(9819 downto 9810) := ADC(11 downto 2);
					when 982 => temp(9829 downto 9820) := ADC(11 downto 2);
					when 983 => temp(9839 downto 9830) := ADC(11 downto 2);
					when 984 => temp(9849 downto 9840) := ADC(11 downto 2);
					when 985 => temp(9859 downto 9850) := ADC(11 downto 2);
					when 986 => temp(9869 downto 9860) := ADC(11 downto 2);
					when 987 => temp(9879 downto 9870) := ADC(11 downto 2);
					when 988 => temp(9889 downto 9880) := ADC(11 downto 2);
					when 989 => temp(9899 downto 9890) := ADC(11 downto 2);
					when 990 => temp(9909 downto 9900) := ADC(11 downto 2);
					when 991 => temp(9919 downto 9910) := ADC(11 downto 2);
					when 992 => temp(9929 downto 9920) := ADC(11 downto 2);
					when 993 => temp(9939 downto 9930) := ADC(11 downto 2);
					when 994 => temp(9949 downto 9940) := ADC(11 downto 2);
					when 995 => temp(9959 downto 9950) := ADC(11 downto 2);
					when 996 => temp(9969 downto 9960) := ADC(11 downto 2);
					when 997 => temp(9979 downto 9970) := ADC(11 downto 2);
					when 998 => temp(9989 downto 9980) := ADC(11 downto 2);
					when 999 => temp(9999 downto 9990) := ADC(11 downto 2);
					when 1000 => temp(10009 downto 10000) := ADC(11 downto 2);
					when 1001 => temp(10019 downto 10010) := ADC(11 downto 2);
					when 1002 => temp(10029 downto 10020) := ADC(11 downto 2);
					when 1003 => temp(10039 downto 10030) := ADC(11 downto 2);
					when 1004 => temp(10049 downto 10040) := ADC(11 downto 2);
					when 1005 => temp(10059 downto 10050) := ADC(11 downto 2);
					when 1006 => temp(10069 downto 10060) := ADC(11 downto 2);
					when 1007 => temp(10079 downto 10070) := ADC(11 downto 2);
					when 1008 => temp(10089 downto 10080) := ADC(11 downto 2);
					when 1009 => temp(10099 downto 10090) := ADC(11 downto 2);
					when 1010 => temp(10109 downto 10100) := ADC(11 downto 2);
					when 1011 => temp(10119 downto 10110) := ADC(11 downto 2);
					when 1012 => temp(10129 downto 10120) := ADC(11 downto 2);
					when 1013 => temp(10139 downto 10130) := ADC(11 downto 2);
					when 1014 => temp(10149 downto 10140) := ADC(11 downto 2);
					when 1015 => temp(10159 downto 10150) := ADC(11 downto 2);
					when 1016 => temp(10169 downto 10160) := ADC(11 downto 2);
					when 1017 => temp(10179 downto 10170) := ADC(11 downto 2);
					when 1018 => temp(10189 downto 10180) := ADC(11 downto 2);
					when 1019 => temp(10199 downto 10190) := ADC(11 downto 2);
					when 1020 => temp(10209 downto 10200) := ADC(11 downto 2);
					when 1021 => temp(10219 downto 10210) := ADC(11 downto 2);
					when 1022 => temp(10229 downto 10220) := ADC(11 downto 2);
					when 1023 => temp(10239 downto 10230) := ADC(11 downto 2);
					when 1024 => temp(10249 downto 10240) := ADC(11 downto 2);
					when 1025 => temp(10259 downto 10250) := ADC(11 downto 2);
					when 1026 => temp(10269 downto 10260) := ADC(11 downto 2);
					when 1027 => temp(10279 downto 10270) := ADC(11 downto 2);
					when 1028 => temp(10289 downto 10280) := ADC(11 downto 2);
					when 1029 => temp(10299 downto 10290) := ADC(11 downto 2);
					when 1030 => temp(10309 downto 10300) := ADC(11 downto 2);
					when 1031 => temp(10319 downto 10310) := ADC(11 downto 2);
					when 1032 => temp(10329 downto 10320) := ADC(11 downto 2);
					when 1033 => temp(10339 downto 10330) := ADC(11 downto 2);
					when 1034 => temp(10349 downto 10340) := ADC(11 downto 2);
					when 1035 => temp(10359 downto 10350) := ADC(11 downto 2);
					when 1036 => temp(10369 downto 10360) := ADC(11 downto 2);
					when 1037 => temp(10379 downto 10370) := ADC(11 downto 2);
					when 1038 => temp(10389 downto 10380) := ADC(11 downto 2);
					when 1039 => temp(10399 downto 10390) := ADC(11 downto 2);
					when 1040 => temp(10409 downto 10400) := ADC(11 downto 2);
					when 1041 => temp(10419 downto 10410) := ADC(11 downto 2);
					when 1042 => temp(10429 downto 10420) := ADC(11 downto 2);
					when 1043 => temp(10439 downto 10430) := ADC(11 downto 2);
					when 1044 => temp(10449 downto 10440) := ADC(11 downto 2);
					when 1045 => temp(10459 downto 10450) := ADC(11 downto 2);
					when 1046 => temp(10469 downto 10460) := ADC(11 downto 2);
					when 1047 => temp(10479 downto 10470) := ADC(11 downto 2);
					when 1048 => temp(10489 downto 10480) := ADC(11 downto 2);
					when 1049 => temp(10499 downto 10490) := ADC(11 downto 2);
					when 1050 => temp(10509 downto 10500) := ADC(11 downto 2);
					when 1051 => temp(10519 downto 10510) := ADC(11 downto 2);
					when 1052 => temp(10529 downto 10520) := ADC(11 downto 2);
					when 1053 => temp(10539 downto 10530) := ADC(11 downto 2);
					when 1054 => temp(10549 downto 10540) := ADC(11 downto 2);
					when 1055 => temp(10559 downto 10550) := ADC(11 downto 2);
					when 1056 => temp(10569 downto 10560) := ADC(11 downto 2);
					when 1057 => temp(10579 downto 10570) := ADC(11 downto 2);
					when 1058 => temp(10589 downto 10580) := ADC(11 downto 2);
					when 1059 => temp(10599 downto 10590) := ADC(11 downto 2);
					when 1060 => temp(10609 downto 10600) := ADC(11 downto 2);
					when 1061 => temp(10619 downto 10610) := ADC(11 downto 2);
					when 1062 => temp(10629 downto 10620) := ADC(11 downto 2);
					when 1063 => temp(10639 downto 10630) := ADC(11 downto 2);
					when 1064 => temp(10649 downto 10640) := ADC(11 downto 2);
					when 1065 => temp(10659 downto 10650) := ADC(11 downto 2);
					when 1066 => temp(10669 downto 10660) := ADC(11 downto 2);
					when 1067 => temp(10679 downto 10670) := ADC(11 downto 2);
					when 1068 => temp(10689 downto 10680) := ADC(11 downto 2);
					when 1069 => temp(10699 downto 10690) := ADC(11 downto 2);
					when 1070 => temp(10709 downto 10700) := ADC(11 downto 2);
					when 1071 => temp(10719 downto 10710) := ADC(11 downto 2);
					when 1072 => temp(10729 downto 10720) := ADC(11 downto 2);
					when 1073 => temp(10739 downto 10730) := ADC(11 downto 2);
					when 1074 => temp(10749 downto 10740) := ADC(11 downto 2);
					when 1075 => temp(10759 downto 10750) := ADC(11 downto 2);
					when 1076 => temp(10769 downto 10760) := ADC(11 downto 2);
					when 1077 => temp(10779 downto 10770) := ADC(11 downto 2);
					when 1078 => temp(10789 downto 10780) := ADC(11 downto 2);
					when 1079 => temp(10799 downto 10790) := ADC(11 downto 2);
					when 1080 => temp(10809 downto 10800) := ADC(11 downto 2);
					when 1081 => temp(10819 downto 10810) := ADC(11 downto 2);
					when 1082 => temp(10829 downto 10820) := ADC(11 downto 2);
					when 1083 => temp(10839 downto 10830) := ADC(11 downto 2);
					when 1084 => temp(10849 downto 10840) := ADC(11 downto 2);
					when 1085 => temp(10859 downto 10850) := ADC(11 downto 2);
					when 1086 => temp(10869 downto 10860) := ADC(11 downto 2);
					when 1087 => temp(10879 downto 10870) := ADC(11 downto 2);
					when 1088 => temp(10889 downto 10880) := ADC(11 downto 2);
					when 1089 => temp(10899 downto 10890) := ADC(11 downto 2);
					when 1090 => temp(10909 downto 10900) := ADC(11 downto 2);
					when 1091 => temp(10919 downto 10910) := ADC(11 downto 2);
					when 1092 => temp(10929 downto 10920) := ADC(11 downto 2);
					when 1093 => temp(10939 downto 10930) := ADC(11 downto 2);
					when 1094 => temp(10949 downto 10940) := ADC(11 downto 2);
					when 1095 => temp(10959 downto 10950) := ADC(11 downto 2);
					when 1096 => temp(10969 downto 10960) := ADC(11 downto 2);
					when 1097 => temp(10979 downto 10970) := ADC(11 downto 2);
					when 1098 => temp(10989 downto 10980) := ADC(11 downto 2);
					when 1099 => temp(10999 downto 10990) := ADC(11 downto 2);
					when 1100 => temp(11009 downto 11000) := ADC(11 downto 2);
					when 1101 => temp(11019 downto 11010) := ADC(11 downto 2);
					when 1102 => temp(11029 downto 11020) := ADC(11 downto 2);
					when 1103 => temp(11039 downto 11030) := ADC(11 downto 2);
					when 1104 => temp(11049 downto 11040) := ADC(11 downto 2);
					when 1105 => temp(11059 downto 11050) := ADC(11 downto 2);
					when 1106 => temp(11069 downto 11060) := ADC(11 downto 2);
					when 1107 => temp(11079 downto 11070) := ADC(11 downto 2);
					when 1108 => temp(11089 downto 11080) := ADC(11 downto 2);
					when 1109 => temp(11099 downto 11090) := ADC(11 downto 2);
					when 1110 => temp(11109 downto 11100) := ADC(11 downto 2);
					when 1111 => temp(11119 downto 11110) := ADC(11 downto 2);
					when 1112 => temp(11129 downto 11120) := ADC(11 downto 2);
					when 1113 => temp(11139 downto 11130) := ADC(11 downto 2);
					when 1114 => temp(11149 downto 11140) := ADC(11 downto 2);
					when 1115 => temp(11159 downto 11150) := ADC(11 downto 2);
					when 1116 => temp(11169 downto 11160) := ADC(11 downto 2);
					when 1117 => temp(11179 downto 11170) := ADC(11 downto 2);
					when 1118 => temp(11189 downto 11180) := ADC(11 downto 2);
					when 1119 => temp(11199 downto 11190) := ADC(11 downto 2);
					when 1120 => temp(11209 downto 11200) := ADC(11 downto 2);
					when 1121 => temp(11219 downto 11210) := ADC(11 downto 2);
					when 1122 => temp(11229 downto 11220) := ADC(11 downto 2);
					when 1123 => temp(11239 downto 11230) := ADC(11 downto 2);
					when 1124 => temp(11249 downto 11240) := ADC(11 downto 2);
					when 1125 => temp(11259 downto 11250) := ADC(11 downto 2);
					when 1126 => temp(11269 downto 11260) := ADC(11 downto 2);
					when 1127 => temp(11279 downto 11270) := ADC(11 downto 2);
					when 1128 => temp(11289 downto 11280) := ADC(11 downto 2);
					when 1129 => temp(11299 downto 11290) := ADC(11 downto 2);
					when 1130 => temp(11309 downto 11300) := ADC(11 downto 2);
					when 1131 => temp(11319 downto 11310) := ADC(11 downto 2);
					when 1132 => temp(11329 downto 11320) := ADC(11 downto 2);
					when 1133 => temp(11339 downto 11330) := ADC(11 downto 2);
					when 1134 => temp(11349 downto 11340) := ADC(11 downto 2);
					when 1135 => temp(11359 downto 11350) := ADC(11 downto 2);
					when 1136 => temp(11369 downto 11360) := ADC(11 downto 2);
					when 1137 => temp(11379 downto 11370) := ADC(11 downto 2);
					when 1138 => temp(11389 downto 11380) := ADC(11 downto 2);
					when 1139 => temp(11399 downto 11390) := ADC(11 downto 2);
					when 1140 => temp(11409 downto 11400) := ADC(11 downto 2);
					when 1141 => temp(11419 downto 11410) := ADC(11 downto 2);
					when 1142 => temp(11429 downto 11420) := ADC(11 downto 2);
					when 1143 => temp(11439 downto 11430) := ADC(11 downto 2);
					when 1144 => temp(11449 downto 11440) := ADC(11 downto 2);
					when 1145 => temp(11459 downto 11450) := ADC(11 downto 2);
					when 1146 => temp(11469 downto 11460) := ADC(11 downto 2);
					when 1147 => temp(11479 downto 11470) := ADC(11 downto 2);
					when 1148 => temp(11489 downto 11480) := ADC(11 downto 2);
					when 1149 => temp(11499 downto 11490) := ADC(11 downto 2);
					when 1150 => temp(11509 downto 11500) := ADC(11 downto 2);
					when 1151 => temp(11519 downto 11510) := ADC(11 downto 2);
					when 1152 => temp(11529 downto 11520) := ADC(11 downto 2);
					when 1153 => temp(11539 downto 11530) := ADC(11 downto 2);
					when 1154 => temp(11549 downto 11540) := ADC(11 downto 2);
					when 1155 => temp(11559 downto 11550) := ADC(11 downto 2);
					when 1156 => temp(11569 downto 11560) := ADC(11 downto 2);
					when 1157 => temp(11579 downto 11570) := ADC(11 downto 2);
					when 1158 => temp(11589 downto 11580) := ADC(11 downto 2);
					when 1159 => temp(11599 downto 11590) := ADC(11 downto 2);
					when 1160 => temp(11609 downto 11600) := ADC(11 downto 2);
					when 1161 => temp(11619 downto 11610) := ADC(11 downto 2);
					when 1162 => temp(11629 downto 11620) := ADC(11 downto 2);
					when 1163 => temp(11639 downto 11630) := ADC(11 downto 2);
					when 1164 => temp(11649 downto 11640) := ADC(11 downto 2);
					when 1165 => temp(11659 downto 11650) := ADC(11 downto 2);
					when 1166 => temp(11669 downto 11660) := ADC(11 downto 2);
					when 1167 => temp(11679 downto 11670) := ADC(11 downto 2);
					when 1168 => temp(11689 downto 11680) := ADC(11 downto 2);
					when 1169 => temp(11699 downto 11690) := ADC(11 downto 2);
					when 1170 => temp(11709 downto 11700) := ADC(11 downto 2);
					when 1171 => temp(11719 downto 11710) := ADC(11 downto 2);
					when 1172 => temp(11729 downto 11720) := ADC(11 downto 2);
					when 1173 => temp(11739 downto 11730) := ADC(11 downto 2);
					when 1174 => temp(11749 downto 11740) := ADC(11 downto 2);
					when 1175 => temp(11759 downto 11750) := ADC(11 downto 2);
					when 1176 => temp(11769 downto 11760) := ADC(11 downto 2);
					when 1177 => temp(11779 downto 11770) := ADC(11 downto 2);
					when 1178 => temp(11789 downto 11780) := ADC(11 downto 2);
					when 1179 => temp(11799 downto 11790) := ADC(11 downto 2);
					when 1180 => temp(11809 downto 11800) := ADC(11 downto 2);
					when 1181 => temp(11819 downto 11810) := ADC(11 downto 2);
					when 1182 => temp(11829 downto 11820) := ADC(11 downto 2);
					when 1183 => temp(11839 downto 11830) := ADC(11 downto 2);
					when 1184 => temp(11849 downto 11840) := ADC(11 downto 2);
					when 1185 => temp(11859 downto 11850) := ADC(11 downto 2);
					when 1186 => temp(11869 downto 11860) := ADC(11 downto 2);
					when 1187 => temp(11879 downto 11870) := ADC(11 downto 2);
					when 1188 => temp(11889 downto 11880) := ADC(11 downto 2);
					when 1189 => temp(11899 downto 11890) := ADC(11 downto 2);
					when 1190 => temp(11909 downto 11900) := ADC(11 downto 2);
					when 1191 => temp(11919 downto 11910) := ADC(11 downto 2);
					when 1192 => temp(11929 downto 11920) := ADC(11 downto 2);
					when 1193 => temp(11939 downto 11930) := ADC(11 downto 2);
					when 1194 => temp(11949 downto 11940) := ADC(11 downto 2);
					when 1195 => temp(11959 downto 11950) := ADC(11 downto 2);
					when 1196 => temp(11969 downto 11960) := ADC(11 downto 2);
					when 1197 => temp(11979 downto 11970) := ADC(11 downto 2);
					when 1198 => temp(11989 downto 11980) := ADC(11 downto 2);
					when 1199 => temp(11999 downto 11990) := ADC(11 downto 2);
					when 1200 => temp(12009 downto 12000) := ADC(11 downto 2);
					when 1201 => temp(12019 downto 12010) := ADC(11 downto 2);
					when 1202 => temp(12029 downto 12020) := ADC(11 downto 2);
					when 1203 => temp(12039 downto 12030) := ADC(11 downto 2);
					when 1204 => temp(12049 downto 12040) := ADC(11 downto 2);
					when 1205 => temp(12059 downto 12050) := ADC(11 downto 2);
					when 1206 => temp(12069 downto 12060) := ADC(11 downto 2);
					when 1207 => temp(12079 downto 12070) := ADC(11 downto 2);
					when 1208 => temp(12089 downto 12080) := ADC(11 downto 2);
					when 1209 => temp(12099 downto 12090) := ADC(11 downto 2);
					when 1210 => temp(12109 downto 12100) := ADC(11 downto 2);
					when 1211 => temp(12119 downto 12110) := ADC(11 downto 2);
					when 1212 => temp(12129 downto 12120) := ADC(11 downto 2);
					when 1213 => temp(12139 downto 12130) := ADC(11 downto 2);
					when 1214 => temp(12149 downto 12140) := ADC(11 downto 2);
					when 1215 => temp(12159 downto 12150) := ADC(11 downto 2);
					when 1216 => temp(12169 downto 12160) := ADC(11 downto 2);
					when 1217 => temp(12179 downto 12170) := ADC(11 downto 2);
					when 1218 => temp(12189 downto 12180) := ADC(11 downto 2);
					when 1219 => temp(12199 downto 12190) := ADC(11 downto 2);
					when 1220 => temp(12209 downto 12200) := ADC(11 downto 2);
					when 1221 => temp(12219 downto 12210) := ADC(11 downto 2);
					when 1222 => temp(12229 downto 12220) := ADC(11 downto 2);
					when 1223 => temp(12239 downto 12230) := ADC(11 downto 2);
					when 1224 => temp(12249 downto 12240) := ADC(11 downto 2);
					when 1225 => temp(12259 downto 12250) := ADC(11 downto 2);
					when 1226 => temp(12269 downto 12260) := ADC(11 downto 2);
					when 1227 => temp(12279 downto 12270) := ADC(11 downto 2);
					when 1228 => temp(12289 downto 12280) := ADC(11 downto 2);
					when 1229 => temp(12299 downto 12290) := ADC(11 downto 2);
					when 1230 => temp(12309 downto 12300) := ADC(11 downto 2);
					when 1231 => temp(12319 downto 12310) := ADC(11 downto 2);
					when 1232 => temp(12329 downto 12320) := ADC(11 downto 2);
					when 1233 => temp(12339 downto 12330) := ADC(11 downto 2);
					when 1234 => temp(12349 downto 12340) := ADC(11 downto 2);
					when 1235 => temp(12359 downto 12350) := ADC(11 downto 2);
					when 1236 => temp(12369 downto 12360) := ADC(11 downto 2);
					when 1237 => temp(12379 downto 12370) := ADC(11 downto 2);
					when 1238 => temp(12389 downto 12380) := ADC(11 downto 2);
					when 1239 => temp(12399 downto 12390) := ADC(11 downto 2);
					when 1240 => temp(12409 downto 12400) := ADC(11 downto 2);
					when 1241 => temp(12419 downto 12410) := ADC(11 downto 2);
					when 1242 => temp(12429 downto 12420) := ADC(11 downto 2);
					when 1243 => temp(12439 downto 12430) := ADC(11 downto 2);
					when 1244 => temp(12449 downto 12440) := ADC(11 downto 2);
					when 1245 => temp(12459 downto 12450) := ADC(11 downto 2);
					when 1246 => temp(12469 downto 12460) := ADC(11 downto 2);
					when 1247 => temp(12479 downto 12470) := ADC(11 downto 2);
					when 1248 => temp(12489 downto 12480) := ADC(11 downto 2);
					when 1249 => temp(12499 downto 12490) := ADC(11 downto 2);
					when 1250 => temp(12509 downto 12500) := ADC(11 downto 2);
					when 1251 => temp(12519 downto 12510) := ADC(11 downto 2);
					when 1252 => temp(12529 downto 12520) := ADC(11 downto 2);
					when 1253 => temp(12539 downto 12530) := ADC(11 downto 2);
					when 1254 => temp(12549 downto 12540) := ADC(11 downto 2);
					when 1255 => temp(12559 downto 12550) := ADC(11 downto 2);
					when 1256 => temp(12569 downto 12560) := ADC(11 downto 2);
					when 1257 => temp(12579 downto 12570) := ADC(11 downto 2);
					when 1258 => temp(12589 downto 12580) := ADC(11 downto 2);
					when 1259 => temp(12599 downto 12590) := ADC(11 downto 2);
					when 1260 => temp(12609 downto 12600) := ADC(11 downto 2);
					when 1261 => temp(12619 downto 12610) := ADC(11 downto 2);
					when 1262 => temp(12629 downto 12620) := ADC(11 downto 2);
					when 1263 => temp(12639 downto 12630) := ADC(11 downto 2);
					when 1264 => temp(12649 downto 12640) := ADC(11 downto 2);
					when 1265 => temp(12659 downto 12650) := ADC(11 downto 2);
					when 1266 => temp(12669 downto 12660) := ADC(11 downto 2);
					when 1267 => temp(12679 downto 12670) := ADC(11 downto 2);
					when 1268 => temp(12689 downto 12680) := ADC(11 downto 2);
					when 1269 => temp(12699 downto 12690) := ADC(11 downto 2);
					when 1270 => temp(12709 downto 12700) := ADC(11 downto 2);
					when 1271 => temp(12719 downto 12710) := ADC(11 downto 2);
					when 1272 => temp(12729 downto 12720) := ADC(11 downto 2);
					when 1273 => temp(12739 downto 12730) := ADC(11 downto 2);
					when 1274 => temp(12749 downto 12740) := ADC(11 downto 2);
					when 1275 => temp(12759 downto 12750) := ADC(11 downto 2);
					when 1276 => temp(12769 downto 12760) := ADC(11 downto 2);
					when 1277 => temp(12779 downto 12770) := ADC(11 downto 2);
					when 1278 => temp(12789 downto 12780) := ADC(11 downto 2);
					when 1279 => temp(12799 downto 12790) := ADC(11 downto 2);
					when 1280 => temp(12809 downto 12800) := ADC(11 downto 2);
					when 1281 => temp(12819 downto 12810) := ADC(11 downto 2);
					when 1282 => temp(12829 downto 12820) := ADC(11 downto 2);
					when 1283 => temp(12839 downto 12830) := ADC(11 downto 2);
					when 1284 => temp(12849 downto 12840) := ADC(11 downto 2);
					when 1285 => temp(12859 downto 12850) := ADC(11 downto 2);
					when 1286 => temp(12869 downto 12860) := ADC(11 downto 2);
					when 1287 => temp(12879 downto 12870) := ADC(11 downto 2);
					when 1288 => temp(12889 downto 12880) := ADC(11 downto 2);
					when 1289 => temp(12899 downto 12890) := ADC(11 downto 2);
					when 1290 => temp(12909 downto 12900) := ADC(11 downto 2);
					when 1291 => temp(12919 downto 12910) := ADC(11 downto 2);
					when 1292 => temp(12929 downto 12920) := ADC(11 downto 2);
					when 1293 => temp(12939 downto 12930) := ADC(11 downto 2);
					when 1294 => temp(12949 downto 12940) := ADC(11 downto 2);
					when 1295 => temp(12959 downto 12950) := ADC(11 downto 2);
					when 1296 => temp(12969 downto 12960) := ADC(11 downto 2);
					when 1297 => temp(12979 downto 12970) := ADC(11 downto 2);
					when 1298 => temp(12989 downto 12980) := ADC(11 downto 2);
					when 1299 => temp(12999 downto 12990) := ADC(11 downto 2);
					when 1300 => temp(13009 downto 13000) := ADC(11 downto 2);
					when 1301 => temp(13019 downto 13010) := ADC(11 downto 2);
					when 1302 => temp(13029 downto 13020) := ADC(11 downto 2);
					when 1303 => temp(13039 downto 13030) := ADC(11 downto 2);
					when 1304 => temp(13049 downto 13040) := ADC(11 downto 2);
					when 1305 => temp(13059 downto 13050) := ADC(11 downto 2);
					when 1306 => temp(13069 downto 13060) := ADC(11 downto 2);
					when 1307 => temp(13079 downto 13070) := ADC(11 downto 2);
					when 1308 => temp(13089 downto 13080) := ADC(11 downto 2);
					when 1309 => temp(13099 downto 13090) := ADC(11 downto 2);
					when 1310 => temp(13109 downto 13100) := ADC(11 downto 2);
					when 1311 => temp(13119 downto 13110) := ADC(11 downto 2);
					when 1312 => temp(13129 downto 13120) := ADC(11 downto 2);
					when 1313 => temp(13139 downto 13130) := ADC(11 downto 2);
					when 1314 => temp(13149 downto 13140) := ADC(11 downto 2);
					when 1315 => temp(13159 downto 13150) := ADC(11 downto 2);
					when 1316 => temp(13169 downto 13160) := ADC(11 downto 2);
					when 1317 => temp(13179 downto 13170) := ADC(11 downto 2);
					when 1318 => temp(13189 downto 13180) := ADC(11 downto 2);
					when 1319 => temp(13199 downto 13190) := ADC(11 downto 2);
					when 1320 => temp(13209 downto 13200) := ADC(11 downto 2);
					when 1321 => temp(13219 downto 13210) := ADC(11 downto 2);
					when 1322 => temp(13229 downto 13220) := ADC(11 downto 2);
					when 1323 => temp(13239 downto 13230) := ADC(11 downto 2);
					when 1324 => temp(13249 downto 13240) := ADC(11 downto 2);
					when 1325 => temp(13259 downto 13250) := ADC(11 downto 2);
					when 1326 => temp(13269 downto 13260) := ADC(11 downto 2);
					when 1327 => temp(13279 downto 13270) := ADC(11 downto 2);
					when 1328 => temp(13289 downto 13280) := ADC(11 downto 2);
					when 1329 => temp(13299 downto 13290) := ADC(11 downto 2);
					when 1330 => temp(13309 downto 13300) := ADC(11 downto 2);
					when 1331 => temp(13319 downto 13310) := ADC(11 downto 2);
					when 1332 => temp(13329 downto 13320) := ADC(11 downto 2);
					when 1333 => temp(13339 downto 13330) := ADC(11 downto 2);
					when 1334 => temp(13349 downto 13340) := ADC(11 downto 2);
					when 1335 => temp(13359 downto 13350) := ADC(11 downto 2);
					when 1336 => temp(13369 downto 13360) := ADC(11 downto 2);
					when 1337 => temp(13379 downto 13370) := ADC(11 downto 2);
					when 1338 => temp(13389 downto 13380) := ADC(11 downto 2);
					when 1339 => temp(13399 downto 13390) := ADC(11 downto 2);
					when 1340 => temp(13409 downto 13400) := ADC(11 downto 2);
					when 1341 => temp(13419 downto 13410) := ADC(11 downto 2);
					when 1342 => temp(13429 downto 13420) := ADC(11 downto 2);
					when 1343 => temp(13439 downto 13430) := ADC(11 downto 2);
					when 1344 => temp(13449 downto 13440) := ADC(11 downto 2);
					when 1345 => temp(13459 downto 13450) := ADC(11 downto 2);
					when 1346 => temp(13469 downto 13460) := ADC(11 downto 2);
					when 1347 => temp(13479 downto 13470) := ADC(11 downto 2);
					when 1348 => temp(13489 downto 13480) := ADC(11 downto 2);
					when 1349 => temp(13499 downto 13490) := ADC(11 downto 2);
					when 1350 => temp(13509 downto 13500) := ADC(11 downto 2);
					when 1351 => temp(13519 downto 13510) := ADC(11 downto 2);
					when 1352 => temp(13529 downto 13520) := ADC(11 downto 2);
					when 1353 => temp(13539 downto 13530) := ADC(11 downto 2);
					when 1354 => temp(13549 downto 13540) := ADC(11 downto 2);
					when 1355 => temp(13559 downto 13550) := ADC(11 downto 2);
					when 1356 => temp(13569 downto 13560) := ADC(11 downto 2);
					when 1357 => temp(13579 downto 13570) := ADC(11 downto 2);
					when 1358 => temp(13589 downto 13580) := ADC(11 downto 2);
					when 1359 => temp(13599 downto 13590) := ADC(11 downto 2);
					when 1360 => temp(13609 downto 13600) := ADC(11 downto 2);
					when 1361 => temp(13619 downto 13610) := ADC(11 downto 2);
					when 1362 => temp(13629 downto 13620) := ADC(11 downto 2);
					when 1363 => temp(13639 downto 13630) := ADC(11 downto 2);
					when 1364 => temp(13649 downto 13640) := ADC(11 downto 2);
					when 1365 => temp(13659 downto 13650) := ADC(11 downto 2);
					when 1366 => temp(13669 downto 13660) := ADC(11 downto 2);
					when 1367 => temp(13679 downto 13670) := ADC(11 downto 2);
					when 1368 => temp(13689 downto 13680) := ADC(11 downto 2);
					when 1369 => temp(13699 downto 13690) := ADC(11 downto 2);
					when 1370 => temp(13709 downto 13700) := ADC(11 downto 2);
					when 1371 => temp(13719 downto 13710) := ADC(11 downto 2);
					when 1372 => temp(13729 downto 13720) := ADC(11 downto 2);
					when 1373 => temp(13739 downto 13730) := ADC(11 downto 2);
					when 1374 => temp(13749 downto 13740) := ADC(11 downto 2);
					when 1375 => temp(13759 downto 13750) := ADC(11 downto 2);
					when 1376 => temp(13769 downto 13760) := ADC(11 downto 2);
					when 1377 => temp(13779 downto 13770) := ADC(11 downto 2);
					when 1378 => temp(13789 downto 13780) := ADC(11 downto 2);
					when 1379 => temp(13799 downto 13790) := ADC(11 downto 2);
					when 1380 => temp(13809 downto 13800) := ADC(11 downto 2);
					when 1381 => temp(13819 downto 13810) := ADC(11 downto 2);
					when 1382 => temp(13829 downto 13820) := ADC(11 downto 2);
					when 1383 => temp(13839 downto 13830) := ADC(11 downto 2);
					when 1384 => temp(13849 downto 13840) := ADC(11 downto 2);
					when 1385 => temp(13859 downto 13850) := ADC(11 downto 2);
					when 1386 => temp(13869 downto 13860) := ADC(11 downto 2);
					when 1387 => temp(13879 downto 13870) := ADC(11 downto 2);
					when 1388 => temp(13889 downto 13880) := ADC(11 downto 2);
					when 1389 => temp(13899 downto 13890) := ADC(11 downto 2);
					when 1390 => temp(13909 downto 13900) := ADC(11 downto 2);
					when 1391 => temp(13919 downto 13910) := ADC(11 downto 2);
					when 1392 => temp(13929 downto 13920) := ADC(11 downto 2);
					when 1393 => temp(13939 downto 13930) := ADC(11 downto 2);
					when 1394 => temp(13949 downto 13940) := ADC(11 downto 2);
					when 1395 => temp(13959 downto 13950) := ADC(11 downto 2);
					when 1396 => temp(13969 downto 13960) := ADC(11 downto 2);
					when 1397 => temp(13979 downto 13970) := ADC(11 downto 2);
					when 1398 => temp(13989 downto 13980) := ADC(11 downto 2);
					when 1399 => temp(13999 downto 13990) := ADC(11 downto 2);
					when 1400 => temp(14009 downto 14000) := ADC(11 downto 2);
					when 1401 => temp(14019 downto 14010) := ADC(11 downto 2);
					when 1402 => temp(14029 downto 14020) := ADC(11 downto 2);
					when 1403 => temp(14039 downto 14030) := ADC(11 downto 2);
					when 1404 => temp(14049 downto 14040) := ADC(11 downto 2);
					when 1405 => temp(14059 downto 14050) := ADC(11 downto 2);
					when 1406 => temp(14069 downto 14060) := ADC(11 downto 2);
					when 1407 => temp(14079 downto 14070) := ADC(11 downto 2);
					when 1408 => temp(14089 downto 14080) := ADC(11 downto 2);
					when 1409 => temp(14099 downto 14090) := ADC(11 downto 2);
					when 1410 => temp(14109 downto 14100) := ADC(11 downto 2);
					when 1411 => temp(14119 downto 14110) := ADC(11 downto 2);
					when 1412 => temp(14129 downto 14120) := ADC(11 downto 2);
					when 1413 => temp(14139 downto 14130) := ADC(11 downto 2);
					when 1414 => temp(14149 downto 14140) := ADC(11 downto 2);
					when 1415 => temp(14159 downto 14150) := ADC(11 downto 2);
					when 1416 => temp(14169 downto 14160) := ADC(11 downto 2);
					when 1417 => temp(14179 downto 14170) := ADC(11 downto 2);
					when 1418 => temp(14189 downto 14180) := ADC(11 downto 2);
					when 1419 => temp(14199 downto 14190) := ADC(11 downto 2);
					when 1420 => temp(14209 downto 14200) := ADC(11 downto 2);
					when 1421 => temp(14219 downto 14210) := ADC(11 downto 2);
					when 1422 => temp(14229 downto 14220) := ADC(11 downto 2);
					when 1423 => temp(14239 downto 14230) := ADC(11 downto 2);
					when 1424 => temp(14249 downto 14240) := ADC(11 downto 2);
					when 1425 => temp(14259 downto 14250) := ADC(11 downto 2);
					when 1426 => temp(14269 downto 14260) := ADC(11 downto 2);
					when 1427 => temp(14279 downto 14270) := ADC(11 downto 2);
					when 1428 => temp(14289 downto 14280) := ADC(11 downto 2);
					when 1429 => temp(14299 downto 14290) := ADC(11 downto 2);
					when 1430 => temp(14309 downto 14300) := ADC(11 downto 2);
					when 1431 => temp(14319 downto 14310) := ADC(11 downto 2);
					when 1432 => temp(14329 downto 14320) := ADC(11 downto 2);
					when 1433 => temp(14339 downto 14330) := ADC(11 downto 2);
					when 1434 => temp(14349 downto 14340) := ADC(11 downto 2);
					when 1435 => temp(14359 downto 14350) := ADC(11 downto 2);
					when 1436 => temp(14369 downto 14360) := ADC(11 downto 2);
					when 1437 => temp(14379 downto 14370) := ADC(11 downto 2);
					when 1438 => temp(14389 downto 14380) := ADC(11 downto 2);
					when 1439 => temp(14399 downto 14390) := ADC(11 downto 2);
					when 1440 => temp(14409 downto 14400) := ADC(11 downto 2);
					when 1441 => temp(14419 downto 14410) := ADC(11 downto 2);
					when 1442 => temp(14429 downto 14420) := ADC(11 downto 2);
					when 1443 => temp(14439 downto 14430) := ADC(11 downto 2);
					when 1444 => temp(14449 downto 14440) := ADC(11 downto 2);
					when 1445 => temp(14459 downto 14450) := ADC(11 downto 2);
					when 1446 => temp(14469 downto 14460) := ADC(11 downto 2);
					when 1447 => temp(14479 downto 14470) := ADC(11 downto 2);
					when 1448 => temp(14489 downto 14480) := ADC(11 downto 2);
					when 1449 => temp(14499 downto 14490) := ADC(11 downto 2);
					when 1450 => temp(14509 downto 14500) := ADC(11 downto 2);
					when 1451 => temp(14519 downto 14510) := ADC(11 downto 2);
					when 1452 => temp(14529 downto 14520) := ADC(11 downto 2);
					when 1453 => temp(14539 downto 14530) := ADC(11 downto 2);
					when 1454 => temp(14549 downto 14540) := ADC(11 downto 2);
					when 1455 => temp(14559 downto 14550) := ADC(11 downto 2);
					when 1456 => temp(14569 downto 14560) := ADC(11 downto 2);
					when 1457 => temp(14579 downto 14570) := ADC(11 downto 2);
					when 1458 => temp(14589 downto 14580) := ADC(11 downto 2);
					when 1459 => temp(14599 downto 14590) := ADC(11 downto 2);
					when 1460 => temp(14609 downto 14600) := ADC(11 downto 2);
					when 1461 => temp(14619 downto 14610) := ADC(11 downto 2);
					when 1462 => temp(14629 downto 14620) := ADC(11 downto 2);
					when 1463 => temp(14639 downto 14630) := ADC(11 downto 2);
					when 1464 => temp(14649 downto 14640) := ADC(11 downto 2);
					when 1465 => temp(14659 downto 14650) := ADC(11 downto 2);
					when 1466 => temp(14669 downto 14660) := ADC(11 downto 2);
					when 1467 => temp(14679 downto 14670) := ADC(11 downto 2);
					when 1468 => temp(14689 downto 14680) := ADC(11 downto 2);
					when 1469 => temp(14699 downto 14690) := ADC(11 downto 2);
					when 1470 => temp(14709 downto 14700) := ADC(11 downto 2);
					when 1471 => temp(14719 downto 14710) := ADC(11 downto 2);
					when 1472 => temp(14729 downto 14720) := ADC(11 downto 2);
					when 1473 => temp(14739 downto 14730) := ADC(11 downto 2);
					when 1474 => temp(14749 downto 14740) := ADC(11 downto 2);
					when 1475 => temp(14759 downto 14750) := ADC(11 downto 2);
					when 1476 => temp(14769 downto 14760) := ADC(11 downto 2);
					when 1477 => temp(14779 downto 14770) := ADC(11 downto 2);
					when 1478 => temp(14789 downto 14780) := ADC(11 downto 2);
					when 1479 => temp(14799 downto 14790) := ADC(11 downto 2);
					when 1480 => temp(14809 downto 14800) := ADC(11 downto 2);
					when 1481 => temp(14819 downto 14810) := ADC(11 downto 2);
					when 1482 => temp(14829 downto 14820) := ADC(11 downto 2);
					when 1483 => temp(14839 downto 14830) := ADC(11 downto 2);
					when 1484 => temp(14849 downto 14840) := ADC(11 downto 2);
					when 1485 => temp(14859 downto 14850) := ADC(11 downto 2);
					when 1486 => temp(14869 downto 14860) := ADC(11 downto 2);
					when 1487 => temp(14879 downto 14870) := ADC(11 downto 2);
					when 1488 => temp(14889 downto 14880) := ADC(11 downto 2);
					when 1489 => temp(14899 downto 14890) := ADC(11 downto 2);
					when 1490 => temp(14909 downto 14900) := ADC(11 downto 2);
					when 1491 => temp(14919 downto 14910) := ADC(11 downto 2);
					when 1492 => temp(14929 downto 14920) := ADC(11 downto 2);
					when 1493 => temp(14939 downto 14930) := ADC(11 downto 2);
					when 1494 => temp(14949 downto 14940) := ADC(11 downto 2);
					when 1495 => temp(14959 downto 14950) := ADC(11 downto 2);
					when 1496 => temp(14969 downto 14960) := ADC(11 downto 2);
					when 1497 => temp(14979 downto 14970) := ADC(11 downto 2);
					when 1498 => temp(14989 downto 14980) := ADC(11 downto 2);
					when 1499 => temp(14999 downto 14990) := ADC(11 downto 2);
					when 1500 => temp(15009 downto 15000) := ADC(11 downto 2);
					when 1501 => temp(15019 downto 15010) := ADC(11 downto 2);
					when 1502 => temp(15029 downto 15020) := ADC(11 downto 2);
					when 1503 => temp(15039 downto 15030) := ADC(11 downto 2);
					when 1504 => temp(15049 downto 15040) := ADC(11 downto 2);
					when 1505 => temp(15059 downto 15050) := ADC(11 downto 2);
					when 1506 => temp(15069 downto 15060) := ADC(11 downto 2);
					when 1507 => temp(15079 downto 15070) := ADC(11 downto 2);
					when 1508 => temp(15089 downto 15080) := ADC(11 downto 2);
					when 1509 => temp(15099 downto 15090) := ADC(11 downto 2);
					when 1510 => temp(15109 downto 15100) := ADC(11 downto 2);
					when 1511 => temp(15119 downto 15110) := ADC(11 downto 2);
					when 1512 => temp(15129 downto 15120) := ADC(11 downto 2);
					when 1513 => temp(15139 downto 15130) := ADC(11 downto 2);
					when 1514 => temp(15149 downto 15140) := ADC(11 downto 2);
					when 1515 => temp(15159 downto 15150) := ADC(11 downto 2);
					when 1516 => temp(15169 downto 15160) := ADC(11 downto 2);
					when 1517 => temp(15179 downto 15170) := ADC(11 downto 2);
					when 1518 => temp(15189 downto 15180) := ADC(11 downto 2);
					when 1519 => temp(15199 downto 15190) := ADC(11 downto 2);
					when 1520 => temp(15209 downto 15200) := ADC(11 downto 2);
					when 1521 => temp(15219 downto 15210) := ADC(11 downto 2);
					when 1522 => temp(15229 downto 15220) := ADC(11 downto 2);
					when 1523 => temp(15239 downto 15230) := ADC(11 downto 2);
					when 1524 => temp(15249 downto 15240) := ADC(11 downto 2);
					when 1525 => temp(15259 downto 15250) := ADC(11 downto 2);
					when 1526 => temp(15269 downto 15260) := ADC(11 downto 2);
					when 1527 => temp(15279 downto 15270) := ADC(11 downto 2);
					when 1528 => temp(15289 downto 15280) := ADC(11 downto 2);
					when 1529 => temp(15299 downto 15290) := ADC(11 downto 2);
					when 1530 => temp(15309 downto 15300) := ADC(11 downto 2);
					when 1531 => temp(15319 downto 15310) := ADC(11 downto 2);
					when 1532 => temp(15329 downto 15320) := ADC(11 downto 2);
					when 1533 => temp(15339 downto 15330) := ADC(11 downto 2);
					when 1534 => temp(15349 downto 15340) := ADC(11 downto 2);
					when 1535 => temp(15359 downto 15350) := ADC(11 downto 2);
					when 1536 => temp(15369 downto 15360) := ADC(11 downto 2);
					when 1537 => temp(15379 downto 15370) := ADC(11 downto 2);
					when 1538 => temp(15389 downto 15380) := ADC(11 downto 2);
					when 1539 => temp(15399 downto 15390) := ADC(11 downto 2);
					when 1540 => temp(15409 downto 15400) := ADC(11 downto 2);
					when 1541 => temp(15419 downto 15410) := ADC(11 downto 2);
					when 1542 => temp(15429 downto 15420) := ADC(11 downto 2);
					when 1543 => temp(15439 downto 15430) := ADC(11 downto 2);
					when 1544 => temp(15449 downto 15440) := ADC(11 downto 2);
					when 1545 => temp(15459 downto 15450) := ADC(11 downto 2);
					when 1546 => temp(15469 downto 15460) := ADC(11 downto 2);
					when 1547 => temp(15479 downto 15470) := ADC(11 downto 2);
					when 1548 => temp(15489 downto 15480) := ADC(11 downto 2);
					when 1549 => temp(15499 downto 15490) := ADC(11 downto 2);
					when 1550 => temp(15509 downto 15500) := ADC(11 downto 2);
					when 1551 => temp(15519 downto 15510) := ADC(11 downto 2);
					when 1552 => temp(15529 downto 15520) := ADC(11 downto 2);
					when 1553 => temp(15539 downto 15530) := ADC(11 downto 2);
					when 1554 => temp(15549 downto 15540) := ADC(11 downto 2);
					when 1555 => temp(15559 downto 15550) := ADC(11 downto 2);
					when 1556 => temp(15569 downto 15560) := ADC(11 downto 2);
					when 1557 => temp(15579 downto 15570) := ADC(11 downto 2);
					when 1558 => temp(15589 downto 15580) := ADC(11 downto 2);
					when 1559 => temp(15599 downto 15590) := ADC(11 downto 2);
					when 1560 => temp(15609 downto 15600) := ADC(11 downto 2);
					when 1561 => temp(15619 downto 15610) := ADC(11 downto 2);
					when 1562 => temp(15629 downto 15620) := ADC(11 downto 2);
					when 1563 => temp(15639 downto 15630) := ADC(11 downto 2);
					when 1564 => temp(15649 downto 15640) := ADC(11 downto 2);
					when 1565 => temp(15659 downto 15650) := ADC(11 downto 2);
					when 1566 => temp(15669 downto 15660) := ADC(11 downto 2);
					when 1567 => temp(15679 downto 15670) := ADC(11 downto 2);
					when 1568 => temp(15689 downto 15680) := ADC(11 downto 2);
					when 1569 => temp(15699 downto 15690) := ADC(11 downto 2);
					when 1570 => temp(15709 downto 15700) := ADC(11 downto 2);
					when 1571 => temp(15719 downto 15710) := ADC(11 downto 2);
					when 1572 => temp(15729 downto 15720) := ADC(11 downto 2);
					when 1573 => temp(15739 downto 15730) := ADC(11 downto 2);
					when 1574 => temp(15749 downto 15740) := ADC(11 downto 2);
					when 1575 => temp(15759 downto 15750) := ADC(11 downto 2);
					when 1576 => temp(15769 downto 15760) := ADC(11 downto 2);
					when 1577 => temp(15779 downto 15770) := ADC(11 downto 2);
					when 1578 => temp(15789 downto 15780) := ADC(11 downto 2);
					when 1579 => temp(15799 downto 15790) := ADC(11 downto 2);
					when 1580 => temp(15809 downto 15800) := ADC(11 downto 2);
					when 1581 => temp(15819 downto 15810) := ADC(11 downto 2);
					when 1582 => temp(15829 downto 15820) := ADC(11 downto 2);
					when 1583 => temp(15839 downto 15830) := ADC(11 downto 2);
					when 1584 => temp(15849 downto 15840) := ADC(11 downto 2);
					when 1585 => temp(15859 downto 15850) := ADC(11 downto 2);
					when 1586 => temp(15869 downto 15860) := ADC(11 downto 2);
					when 1587 => temp(15879 downto 15870) := ADC(11 downto 2);
					when 1588 => temp(15889 downto 15880) := ADC(11 downto 2);
					when 1589 => temp(15899 downto 15890) := ADC(11 downto 2);
					when 1590 => temp(15909 downto 15900) := ADC(11 downto 2);
					when 1591 => temp(15919 downto 15910) := ADC(11 downto 2);
					when 1592 => temp(15929 downto 15920) := ADC(11 downto 2);
					when 1593 => temp(15939 downto 15930) := ADC(11 downto 2);
					when 1594 => temp(15949 downto 15940) := ADC(11 downto 2);
					when 1595 => temp(15959 downto 15950) := ADC(11 downto 2);
					when 1596 => temp(15969 downto 15960) := ADC(11 downto 2);
					when 1597 => temp(15979 downto 15970) := ADC(11 downto 2);
					when 1598 => temp(15989 downto 15980) := ADC(11 downto 2);
					when 1599 => temp(15999 downto 15990) := ADC(11 downto 2);
					when 1600 => temp(16009 downto 16000) := ADC(11 downto 2);
					when 1601 => temp(16019 downto 16010) := ADC(11 downto 2);
					when 1602 => temp(16029 downto 16020) := ADC(11 downto 2);
					when 1603 => temp(16039 downto 16030) := ADC(11 downto 2);
					when 1604 => temp(16049 downto 16040) := ADC(11 downto 2);
					when 1605 => temp(16059 downto 16050) := ADC(11 downto 2);
					when 1606 => temp(16069 downto 16060) := ADC(11 downto 2);
					when 1607 => temp(16079 downto 16070) := ADC(11 downto 2);
					when 1608 => temp(16089 downto 16080) := ADC(11 downto 2);
					when 1609 => temp(16099 downto 16090) := ADC(11 downto 2);
					when 1610 => temp(16109 downto 16100) := ADC(11 downto 2);
					when 1611 => temp(16119 downto 16110) := ADC(11 downto 2);
					when 1612 => temp(16129 downto 16120) := ADC(11 downto 2);
					when 1613 => temp(16139 downto 16130) := ADC(11 downto 2);
					when 1614 => temp(16149 downto 16140) := ADC(11 downto 2);
					when 1615 => temp(16159 downto 16150) := ADC(11 downto 2);
					when 1616 => temp(16169 downto 16160) := ADC(11 downto 2);
					when 1617 => temp(16179 downto 16170) := ADC(11 downto 2);
					when 1618 => temp(16189 downto 16180) := ADC(11 downto 2);
					when 1619 => temp(16199 downto 16190) := ADC(11 downto 2);
					when 1620 => temp(16209 downto 16200) := ADC(11 downto 2);
					when 1621 => temp(16219 downto 16210) := ADC(11 downto 2);
					when 1622 => temp(16229 downto 16220) := ADC(11 downto 2);
					when 1623 => temp(16239 downto 16230) := ADC(11 downto 2);
					when 1624 => temp(16249 downto 16240) := ADC(11 downto 2);
					when 1625 => temp(16259 downto 16250) := ADC(11 downto 2);
					when 1626 => temp(16269 downto 16260) := ADC(11 downto 2);
					when 1627 => temp(16279 downto 16270) := ADC(11 downto 2);
					when 1628 => temp(16289 downto 16280) := ADC(11 downto 2);
					when 1629 => temp(16299 downto 16290) := ADC(11 downto 2);
					when 1630 => temp(16309 downto 16300) := ADC(11 downto 2);
					when 1631 => temp(16319 downto 16310) := ADC(11 downto 2);
					when 1632 => temp(16329 downto 16320) := ADC(11 downto 2);
					when 1633 => temp(16339 downto 16330) := ADC(11 downto 2);
					when 1634 => temp(16349 downto 16340) := ADC(11 downto 2);
					when 1635 => temp(16359 downto 16350) := ADC(11 downto 2);
					when 1636 => temp(16369 downto 16360) := ADC(11 downto 2);
					when 1637 => temp(16379 downto 16370) := ADC(11 downto 2);
					when 1638 => temp(16389 downto 16380) := ADC(11 downto 2);
					when 1639 => temp(16399 downto 16390) := ADC(11 downto 2);
					when 1640 => temp(16409 downto 16400) := ADC(11 downto 2);
					when 1641 => temp(16419 downto 16410) := ADC(11 downto 2);
					when 1642 => temp(16429 downto 16420) := ADC(11 downto 2);
					when 1643 => temp(16439 downto 16430) := ADC(11 downto 2);
					when 1644 => temp(16449 downto 16440) := ADC(11 downto 2);
					when 1645 => temp(16459 downto 16450) := ADC(11 downto 2);
					when 1646 => temp(16469 downto 16460) := ADC(11 downto 2);
					when 1647 => temp(16479 downto 16470) := ADC(11 downto 2);
					when 1648 => temp(16489 downto 16480) := ADC(11 downto 2);
					when 1649 => temp(16499 downto 16490) := ADC(11 downto 2);
					when 1650 => temp(16509 downto 16500) := ADC(11 downto 2);
					when 1651 => temp(16519 downto 16510) := ADC(11 downto 2);
					when 1652 => temp(16529 downto 16520) := ADC(11 downto 2);
					when 1653 => temp(16539 downto 16530) := ADC(11 downto 2);
					when 1654 => temp(16549 downto 16540) := ADC(11 downto 2);
					when 1655 => temp(16559 downto 16550) := ADC(11 downto 2);
					when 1656 => temp(16569 downto 16560) := ADC(11 downto 2);
					when 1657 => temp(16579 downto 16570) := ADC(11 downto 2);
					when 1658 => temp(16589 downto 16580) := ADC(11 downto 2);
					when 1659 => temp(16599 downto 16590) := ADC(11 downto 2);
					when 1660 => temp(16609 downto 16600) := ADC(11 downto 2);
					when 1661 => temp(16619 downto 16610) := ADC(11 downto 2);
					when 1662 => temp(16629 downto 16620) := ADC(11 downto 2);
					when 1663 => temp(16639 downto 16630) := ADC(11 downto 2);
					when 1664 => temp(16649 downto 16640) := ADC(11 downto 2);
					when 1665 => temp(16659 downto 16650) := ADC(11 downto 2);
					when 1666 => temp(16669 downto 16660) := ADC(11 downto 2);
					when 1667 => temp(16679 downto 16670) := ADC(11 downto 2);
					when 1668 => temp(16689 downto 16680) := ADC(11 downto 2);
					when 1669 => temp(16699 downto 16690) := ADC(11 downto 2);
					when 1670 => temp(16709 downto 16700) := ADC(11 downto 2);
					when 1671 => temp(16719 downto 16710) := ADC(11 downto 2);
					when 1672 => temp(16729 downto 16720) := ADC(11 downto 2);
					when 1673 => temp(16739 downto 16730) := ADC(11 downto 2);
					when 1674 => temp(16749 downto 16740) := ADC(11 downto 2);
					when 1675 => temp(16759 downto 16750) := ADC(11 downto 2);
					when 1676 => temp(16769 downto 16760) := ADC(11 downto 2);
					when 1677 => temp(16779 downto 16770) := ADC(11 downto 2);
					when 1678 => temp(16789 downto 16780) := ADC(11 downto 2);
					when 1679 => temp(16799 downto 16790) := ADC(11 downto 2);
					when 1680 => temp(16809 downto 16800) := ADC(11 downto 2);
					when 1681 => temp(16819 downto 16810) := ADC(11 downto 2);
					when 1682 => temp(16829 downto 16820) := ADC(11 downto 2);
					when 1683 => temp(16839 downto 16830) := ADC(11 downto 2);
					when 1684 => temp(16849 downto 16840) := ADC(11 downto 2);
					when 1685 => temp(16859 downto 16850) := ADC(11 downto 2);
					when 1686 => temp(16869 downto 16860) := ADC(11 downto 2);
					when 1687 => temp(16879 downto 16870) := ADC(11 downto 2);
					when 1688 => temp(16889 downto 16880) := ADC(11 downto 2);
					when 1689 => temp(16899 downto 16890) := ADC(11 downto 2);
					when 1690 => temp(16909 downto 16900) := ADC(11 downto 2);
					when 1691 => temp(16919 downto 16910) := ADC(11 downto 2);
					when 1692 => temp(16929 downto 16920) := ADC(11 downto 2);
					when 1693 => temp(16939 downto 16930) := ADC(11 downto 2);
					when 1694 => temp(16949 downto 16940) := ADC(11 downto 2);
					when 1695 => temp(16959 downto 16950) := ADC(11 downto 2);
					when 1696 => temp(16969 downto 16960) := ADC(11 downto 2);
					when 1697 => temp(16979 downto 16970) := ADC(11 downto 2);
					when 1698 => temp(16989 downto 16980) := ADC(11 downto 2);
					when 1699 => temp(16999 downto 16990) := ADC(11 downto 2);
					when 1700 => temp(17009 downto 17000) := ADC(11 downto 2);
					when 1701 => temp(17019 downto 17010) := ADC(11 downto 2);
					when 1702 => temp(17029 downto 17020) := ADC(11 downto 2);
					when 1703 => temp(17039 downto 17030) := ADC(11 downto 2);
					when 1704 => temp(17049 downto 17040) := ADC(11 downto 2);
					when 1705 => temp(17059 downto 17050) := ADC(11 downto 2);
					when 1706 => temp(17069 downto 17060) := ADC(11 downto 2);
					when 1707 => temp(17079 downto 17070) := ADC(11 downto 2);
					when 1708 => temp(17089 downto 17080) := ADC(11 downto 2);
					when 1709 => temp(17099 downto 17090) := ADC(11 downto 2);
					when 1710 => temp(17109 downto 17100) := ADC(11 downto 2);
					when 1711 => temp(17119 downto 17110) := ADC(11 downto 2);
					when 1712 => temp(17129 downto 17120) := ADC(11 downto 2);
					when 1713 => temp(17139 downto 17130) := ADC(11 downto 2);
					when 1714 => temp(17149 downto 17140) := ADC(11 downto 2);
					when 1715 => temp(17159 downto 17150) := ADC(11 downto 2);
					when 1716 => temp(17169 downto 17160) := ADC(11 downto 2);
					when 1717 => temp(17179 downto 17170) := ADC(11 downto 2);
					when 1718 => temp(17189 downto 17180) := ADC(11 downto 2);
					when 1719 => temp(17199 downto 17190) := ADC(11 downto 2);
					when 1720 => temp(17209 downto 17200) := ADC(11 downto 2);
					when 1721 => temp(17219 downto 17210) := ADC(11 downto 2);
					when 1722 => temp(17229 downto 17220) := ADC(11 downto 2);
					when 1723 => temp(17239 downto 17230) := ADC(11 downto 2);
					when 1724 => temp(17249 downto 17240) := ADC(11 downto 2);
					when 1725 => temp(17259 downto 17250) := ADC(11 downto 2);
					when 1726 => temp(17269 downto 17260) := ADC(11 downto 2);
					when 1727 => temp(17279 downto 17270) := ADC(11 downto 2);
					when 1728 => temp(17289 downto 17280) := ADC(11 downto 2);
					when 1729 => temp(17299 downto 17290) := ADC(11 downto 2);
					when 1730 => temp(17309 downto 17300) := ADC(11 downto 2);
					when 1731 => temp(17319 downto 17310) := ADC(11 downto 2);
					when 1732 => temp(17329 downto 17320) := ADC(11 downto 2);
					when 1733 => temp(17339 downto 17330) := ADC(11 downto 2);
					when 1734 => temp(17349 downto 17340) := ADC(11 downto 2);
					when 1735 => temp(17359 downto 17350) := ADC(11 downto 2);
					when 1736 => temp(17369 downto 17360) := ADC(11 downto 2);
					when 1737 => temp(17379 downto 17370) := ADC(11 downto 2);
					when 1738 => temp(17389 downto 17380) := ADC(11 downto 2);
					when 1739 => temp(17399 downto 17390) := ADC(11 downto 2);
					when 1740 => temp(17409 downto 17400) := ADC(11 downto 2);
					when 1741 => temp(17419 downto 17410) := ADC(11 downto 2);
					when 1742 => temp(17429 downto 17420) := ADC(11 downto 2);
					when 1743 => temp(17439 downto 17430) := ADC(11 downto 2);
					when 1744 => temp(17449 downto 17440) := ADC(11 downto 2);
					when 1745 => temp(17459 downto 17450) := ADC(11 downto 2);
					when 1746 => temp(17469 downto 17460) := ADC(11 downto 2);
					when 1747 => temp(17479 downto 17470) := ADC(11 downto 2);
					when 1748 => temp(17489 downto 17480) := ADC(11 downto 2);
					when 1749 => temp(17499 downto 17490) := ADC(11 downto 2);
					when 1750 => temp(17509 downto 17500) := ADC(11 downto 2);
					when 1751 => temp(17519 downto 17510) := ADC(11 downto 2);
					when 1752 => temp(17529 downto 17520) := ADC(11 downto 2);
					when 1753 => temp(17539 downto 17530) := ADC(11 downto 2);
					when 1754 => temp(17549 downto 17540) := ADC(11 downto 2);
					when 1755 => temp(17559 downto 17550) := ADC(11 downto 2);
					when 1756 => temp(17569 downto 17560) := ADC(11 downto 2);
					when 1757 => temp(17579 downto 17570) := ADC(11 downto 2);
					when 1758 => temp(17589 downto 17580) := ADC(11 downto 2);
					when 1759 => temp(17599 downto 17590) := ADC(11 downto 2);
					when 1760 => temp(17609 downto 17600) := ADC(11 downto 2);
					when 1761 => temp(17619 downto 17610) := ADC(11 downto 2);
					when 1762 => temp(17629 downto 17620) := ADC(11 downto 2);
					when 1763 => temp(17639 downto 17630) := ADC(11 downto 2);
					when 1764 => temp(17649 downto 17640) := ADC(11 downto 2);
					when 1765 => temp(17659 downto 17650) := ADC(11 downto 2);
					when 1766 => temp(17669 downto 17660) := ADC(11 downto 2);
					when 1767 => temp(17679 downto 17670) := ADC(11 downto 2);
					when 1768 => temp(17689 downto 17680) := ADC(11 downto 2);
					when 1769 => temp(17699 downto 17690) := ADC(11 downto 2);
					when 1770 => temp(17709 downto 17700) := ADC(11 downto 2);
					when 1771 => temp(17719 downto 17710) := ADC(11 downto 2);
					when 1772 => temp(17729 downto 17720) := ADC(11 downto 2);
					when 1773 => temp(17739 downto 17730) := ADC(11 downto 2);
					when 1774 => temp(17749 downto 17740) := ADC(11 downto 2);
					when 1775 => temp(17759 downto 17750) := ADC(11 downto 2);
					when 1776 => temp(17769 downto 17760) := ADC(11 downto 2);
					when 1777 => temp(17779 downto 17770) := ADC(11 downto 2);
					when 1778 => temp(17789 downto 17780) := ADC(11 downto 2);
					when 1779 => temp(17799 downto 17790) := ADC(11 downto 2);
					when 1780 => temp(17809 downto 17800) := ADC(11 downto 2);
					when 1781 => temp(17819 downto 17810) := ADC(11 downto 2);
					when 1782 => temp(17829 downto 17820) := ADC(11 downto 2);
					when 1783 => temp(17839 downto 17830) := ADC(11 downto 2);
					when 1784 => temp(17849 downto 17840) := ADC(11 downto 2);
					when 1785 => temp(17859 downto 17850) := ADC(11 downto 2);
					when 1786 => temp(17869 downto 17860) := ADC(11 downto 2);
					when 1787 => temp(17879 downto 17870) := ADC(11 downto 2);
					when 1788 => temp(17889 downto 17880) := ADC(11 downto 2);
					when 1789 => temp(17899 downto 17890) := ADC(11 downto 2);
					when 1790 => temp(17909 downto 17900) := ADC(11 downto 2);
					when 1791 => temp(17919 downto 17910) := ADC(11 downto 2);
					when 1792 => temp(17929 downto 17920) := ADC(11 downto 2);
					when 1793 => temp(17939 downto 17930) := ADC(11 downto 2);
					when 1794 => temp(17949 downto 17940) := ADC(11 downto 2);
					when 1795 => temp(17959 downto 17950) := ADC(11 downto 2);
					when 1796 => temp(17969 downto 17960) := ADC(11 downto 2);
					when 1797 => temp(17979 downto 17970) := ADC(11 downto 2);
					when 1798 => temp(17989 downto 17980) := ADC(11 downto 2);
					when 1799 => temp(17999 downto 17990) := ADC(11 downto 2);
					when 1800 => temp(18009 downto 18000) := ADC(11 downto 2);
					when 1801 => temp(18019 downto 18010) := ADC(11 downto 2);
					when 1802 => temp(18029 downto 18020) := ADC(11 downto 2);
					when 1803 => temp(18039 downto 18030) := ADC(11 downto 2);
					when 1804 => temp(18049 downto 18040) := ADC(11 downto 2);
					when 1805 => temp(18059 downto 18050) := ADC(11 downto 2);
					when 1806 => temp(18069 downto 18060) := ADC(11 downto 2);
					when 1807 => temp(18079 downto 18070) := ADC(11 downto 2);
					when 1808 => temp(18089 downto 18080) := ADC(11 downto 2);
					when 1809 => temp(18099 downto 18090) := ADC(11 downto 2);
					when 1810 => temp(18109 downto 18100) := ADC(11 downto 2);
					when 1811 => temp(18119 downto 18110) := ADC(11 downto 2);
					when 1812 => temp(18129 downto 18120) := ADC(11 downto 2);
					when 1813 => temp(18139 downto 18130) := ADC(11 downto 2);
					when 1814 => temp(18149 downto 18140) := ADC(11 downto 2);
					when 1815 => temp(18159 downto 18150) := ADC(11 downto 2);
					when 1816 => temp(18169 downto 18160) := ADC(11 downto 2);
					when 1817 => temp(18179 downto 18170) := ADC(11 downto 2);
					when 1818 => temp(18189 downto 18180) := ADC(11 downto 2);
					when 1819 => temp(18199 downto 18190) := ADC(11 downto 2);
					when 1820 => temp(18209 downto 18200) := ADC(11 downto 2);
					when 1821 => temp(18219 downto 18210) := ADC(11 downto 2);
					when 1822 => temp(18229 downto 18220) := ADC(11 downto 2);
					when 1823 => temp(18239 downto 18230) := ADC(11 downto 2);
					when 1824 => temp(18249 downto 18240) := ADC(11 downto 2);
					when 1825 => temp(18259 downto 18250) := ADC(11 downto 2);
					when 1826 => temp(18269 downto 18260) := ADC(11 downto 2);
					when 1827 => temp(18279 downto 18270) := ADC(11 downto 2);
					when 1828 => temp(18289 downto 18280) := ADC(11 downto 2);
					when 1829 => temp(18299 downto 18290) := ADC(11 downto 2);
					when 1830 => temp(18309 downto 18300) := ADC(11 downto 2);
					when 1831 => temp(18319 downto 18310) := ADC(11 downto 2);
					when 1832 => temp(18329 downto 18320) := ADC(11 downto 2);
					when 1833 => temp(18339 downto 18330) := ADC(11 downto 2);
					when 1834 => temp(18349 downto 18340) := ADC(11 downto 2);
					when 1835 => temp(18359 downto 18350) := ADC(11 downto 2);
					when 1836 => temp(18369 downto 18360) := ADC(11 downto 2);
					when 1837 => temp(18379 downto 18370) := ADC(11 downto 2);
					when 1838 => temp(18389 downto 18380) := ADC(11 downto 2);
					when 1839 => temp(18399 downto 18390) := ADC(11 downto 2);
					when 1840 => temp(18409 downto 18400) := ADC(11 downto 2);
					when 1841 => temp(18419 downto 18410) := ADC(11 downto 2);
					when 1842 => temp(18429 downto 18420) := ADC(11 downto 2);
					when 1843 => temp(18439 downto 18430) := ADC(11 downto 2);
					when 1844 => temp(18449 downto 18440) := ADC(11 downto 2);
					when 1845 => temp(18459 downto 18450) := ADC(11 downto 2);
					when 1846 => temp(18469 downto 18460) := ADC(11 downto 2);
					when 1847 => temp(18479 downto 18470) := ADC(11 downto 2);
					when 1848 => temp(18489 downto 18480) := ADC(11 downto 2);
					when 1849 => temp(18499 downto 18490) := ADC(11 downto 2);
					when 1850 => temp(18509 downto 18500) := ADC(11 downto 2);
					when 1851 => temp(18519 downto 18510) := ADC(11 downto 2);
					when 1852 => temp(18529 downto 18520) := ADC(11 downto 2);
					when 1853 => temp(18539 downto 18530) := ADC(11 downto 2);
					when 1854 => temp(18549 downto 18540) := ADC(11 downto 2);
					when 1855 => temp(18559 downto 18550) := ADC(11 downto 2);
					when 1856 => temp(18569 downto 18560) := ADC(11 downto 2);
					when 1857 => temp(18579 downto 18570) := ADC(11 downto 2);
					when 1858 => temp(18589 downto 18580) := ADC(11 downto 2);
					when 1859 => temp(18599 downto 18590) := ADC(11 downto 2);
					when 1860 => temp(18609 downto 18600) := ADC(11 downto 2);
					when 1861 => temp(18619 downto 18610) := ADC(11 downto 2);
					when 1862 => temp(18629 downto 18620) := ADC(11 downto 2);
					when 1863 => temp(18639 downto 18630) := ADC(11 downto 2);
					when 1864 => temp(18649 downto 18640) := ADC(11 downto 2);
					when 1865 => temp(18659 downto 18650) := ADC(11 downto 2);
					when 1866 => temp(18669 downto 18660) := ADC(11 downto 2);
					when 1867 => temp(18679 downto 18670) := ADC(11 downto 2);
					when 1868 => temp(18689 downto 18680) := ADC(11 downto 2);
					when 1869 => temp(18699 downto 18690) := ADC(11 downto 2);
					when 1870 => temp(18709 downto 18700) := ADC(11 downto 2);
					when 1871 => temp(18719 downto 18710) := ADC(11 downto 2);
					when 1872 => temp(18729 downto 18720) := ADC(11 downto 2);
					when 1873 => temp(18739 downto 18730) := ADC(11 downto 2);
					when 1874 => temp(18749 downto 18740) := ADC(11 downto 2);
					when 1875 => temp(18759 downto 18750) := ADC(11 downto 2);
					when 1876 => temp(18769 downto 18760) := ADC(11 downto 2);
					when 1877 => temp(18779 downto 18770) := ADC(11 downto 2);
					when 1878 => temp(18789 downto 18780) := ADC(11 downto 2);
					when 1879 => temp(18799 downto 18790) := ADC(11 downto 2);
					when 1880 => temp(18809 downto 18800) := ADC(11 downto 2);
					when 1881 => temp(18819 downto 18810) := ADC(11 downto 2);
					when 1882 => temp(18829 downto 18820) := ADC(11 downto 2);
					when 1883 => temp(18839 downto 18830) := ADC(11 downto 2);
					when 1884 => temp(18849 downto 18840) := ADC(11 downto 2);
					when 1885 => temp(18859 downto 18850) := ADC(11 downto 2);
					when 1886 => temp(18869 downto 18860) := ADC(11 downto 2);
					when 1887 => temp(18879 downto 18870) := ADC(11 downto 2);
					when 1888 => temp(18889 downto 18880) := ADC(11 downto 2);
					when 1889 => temp(18899 downto 18890) := ADC(11 downto 2);
					when 1890 => temp(18909 downto 18900) := ADC(11 downto 2);
					when 1891 => temp(18919 downto 18910) := ADC(11 downto 2);
					when 1892 => temp(18929 downto 18920) := ADC(11 downto 2);
					when 1893 => temp(18939 downto 18930) := ADC(11 downto 2);
					when 1894 => temp(18949 downto 18940) := ADC(11 downto 2);
					when 1895 => temp(18959 downto 18950) := ADC(11 downto 2);
					when 1896 => temp(18969 downto 18960) := ADC(11 downto 2);
					when 1897 => temp(18979 downto 18970) := ADC(11 downto 2);
					when 1898 => temp(18989 downto 18980) := ADC(11 downto 2);
					when 1899 => temp(18999 downto 18990) := ADC(11 downto 2);
					when 1900 => temp(19009 downto 19000) := ADC(11 downto 2);
					when 1901 => temp(19019 downto 19010) := ADC(11 downto 2);
					when 1902 => temp(19029 downto 19020) := ADC(11 downto 2);
					when 1903 => temp(19039 downto 19030) := ADC(11 downto 2);
					when 1904 => temp(19049 downto 19040) := ADC(11 downto 2);
					when 1905 => temp(19059 downto 19050) := ADC(11 downto 2);
					when 1906 => temp(19069 downto 19060) := ADC(11 downto 2);
					when 1907 => temp(19079 downto 19070) := ADC(11 downto 2);
					when 1908 => temp(19089 downto 19080) := ADC(11 downto 2);
					when 1909 => temp(19099 downto 19090) := ADC(11 downto 2);
					when 1910 => temp(19109 downto 19100) := ADC(11 downto 2);
					when 1911 => temp(19119 downto 19110) := ADC(11 downto 2);
					when 1912 => temp(19129 downto 19120) := ADC(11 downto 2);
					when 1913 => temp(19139 downto 19130) := ADC(11 downto 2);
					when 1914 => temp(19149 downto 19140) := ADC(11 downto 2);
					when 1915 => temp(19159 downto 19150) := ADC(11 downto 2);
					when 1916 => temp(19169 downto 19160) := ADC(11 downto 2);
					when 1917 => temp(19179 downto 19170) := ADC(11 downto 2);
					when 1918 => temp(19189 downto 19180) := ADC(11 downto 2);
					when 1919 => temp(19199 downto 19190) := ADC(11 downto 2);
					when 1920 => temp(19209 downto 19200) := ADC(11 downto 2);
					when 1921 => temp(19219 downto 19210) := ADC(11 downto 2);
					when 1922 => temp(19229 downto 19220) := ADC(11 downto 2);
					when 1923 => temp(19239 downto 19230) := ADC(11 downto 2);
					when 1924 => temp(19249 downto 19240) := ADC(11 downto 2);
					when 1925 => temp(19259 downto 19250) := ADC(11 downto 2);
					when 1926 => temp(19269 downto 19260) := ADC(11 downto 2);
					when 1927 => temp(19279 downto 19270) := ADC(11 downto 2);
					when 1928 => temp(19289 downto 19280) := ADC(11 downto 2);
					when 1929 => temp(19299 downto 19290) := ADC(11 downto 2);
					when 1930 => temp(19309 downto 19300) := ADC(11 downto 2);
					when 1931 => temp(19319 downto 19310) := ADC(11 downto 2);
					when 1932 => temp(19329 downto 19320) := ADC(11 downto 2);
					when 1933 => temp(19339 downto 19330) := ADC(11 downto 2);
					when 1934 => temp(19349 downto 19340) := ADC(11 downto 2);
					when 1935 => temp(19359 downto 19350) := ADC(11 downto 2);
					when 1936 => temp(19369 downto 19360) := ADC(11 downto 2);
					when 1937 => temp(19379 downto 19370) := ADC(11 downto 2);
					when 1938 => temp(19389 downto 19380) := ADC(11 downto 2);
					when 1939 => temp(19399 downto 19390) := ADC(11 downto 2);
					when 1940 => temp(19409 downto 19400) := ADC(11 downto 2);
					when 1941 => temp(19419 downto 19410) := ADC(11 downto 2);
					when 1942 => temp(19429 downto 19420) := ADC(11 downto 2);
					when 1943 => temp(19439 downto 19430) := ADC(11 downto 2);
					when 1944 => temp(19449 downto 19440) := ADC(11 downto 2);
					when 1945 => temp(19459 downto 19450) := ADC(11 downto 2);
					when 1946 => temp(19469 downto 19460) := ADC(11 downto 2);
					when 1947 => temp(19479 downto 19470) := ADC(11 downto 2);
					when 1948 => temp(19489 downto 19480) := ADC(11 downto 2);
					when 1949 => temp(19499 downto 19490) := ADC(11 downto 2);
					when 1950 => temp(19509 downto 19500) := ADC(11 downto 2);
					when 1951 => temp(19519 downto 19510) := ADC(11 downto 2);
					when 1952 => temp(19529 downto 19520) := ADC(11 downto 2);
					when 1953 => temp(19539 downto 19530) := ADC(11 downto 2);
					when 1954 => temp(19549 downto 19540) := ADC(11 downto 2);
					when 1955 => temp(19559 downto 19550) := ADC(11 downto 2);
					when 1956 => temp(19569 downto 19560) := ADC(11 downto 2);
					when 1957 => temp(19579 downto 19570) := ADC(11 downto 2);
					when 1958 => temp(19589 downto 19580) := ADC(11 downto 2);
					when 1959 => temp(19599 downto 19590) := ADC(11 downto 2);
					when 1960 => temp(19609 downto 19600) := ADC(11 downto 2);
					when 1961 => temp(19619 downto 19610) := ADC(11 downto 2);
					when 1962 => temp(19629 downto 19620) := ADC(11 downto 2);
					when 1963 => temp(19639 downto 19630) := ADC(11 downto 2);
					when 1964 => temp(19649 downto 19640) := ADC(11 downto 2);
					when 1965 => temp(19659 downto 19650) := ADC(11 downto 2);
					when 1966 => temp(19669 downto 19660) := ADC(11 downto 2);
					when 1967 => temp(19679 downto 19670) := ADC(11 downto 2);
					when 1968 => temp(19689 downto 19680) := ADC(11 downto 2);
					when 1969 => temp(19699 downto 19690) := ADC(11 downto 2);
					when 1970 => temp(19709 downto 19700) := ADC(11 downto 2);
					when 1971 => temp(19719 downto 19710) := ADC(11 downto 2);
					when 1972 => temp(19729 downto 19720) := ADC(11 downto 2);
					when 1973 => temp(19739 downto 19730) := ADC(11 downto 2);
					when 1974 => temp(19749 downto 19740) := ADC(11 downto 2);
					when 1975 => temp(19759 downto 19750) := ADC(11 downto 2);
					when 1976 => temp(19769 downto 19760) := ADC(11 downto 2);
					when 1977 => temp(19779 downto 19770) := ADC(11 downto 2);
					when 1978 => temp(19789 downto 19780) := ADC(11 downto 2);
					when 1979 => temp(19799 downto 19790) := ADC(11 downto 2);
					when 1980 => temp(19809 downto 19800) := ADC(11 downto 2);
					when 1981 => temp(19819 downto 19810) := ADC(11 downto 2);
					when 1982 => temp(19829 downto 19820) := ADC(11 downto 2);
					when 1983 => temp(19839 downto 19830) := ADC(11 downto 2);
					when 1984 => temp(19849 downto 19840) := ADC(11 downto 2);
					when 1985 => temp(19859 downto 19850) := ADC(11 downto 2);
					when 1986 => temp(19869 downto 19860) := ADC(11 downto 2);
					when 1987 => temp(19879 downto 19870) := ADC(11 downto 2);
					when 1988 => temp(19889 downto 19880) := ADC(11 downto 2);
					when 1989 => temp(19899 downto 19890) := ADC(11 downto 2);
					when 1990 => temp(19909 downto 19900) := ADC(11 downto 2);
					when 1991 => temp(19919 downto 19910) := ADC(11 downto 2);
					when 1992 => temp(19929 downto 19920) := ADC(11 downto 2);
					when 1993 => temp(19939 downto 19930) := ADC(11 downto 2);
					when 1994 => temp(19949 downto 19940) := ADC(11 downto 2);
					when 1995 => temp(19959 downto 19950) := ADC(11 downto 2);
					when 1996 => temp(19969 downto 19960) := ADC(11 downto 2);
					when 1997 => temp(19979 downto 19970) := ADC(11 downto 2);
					when 1998 => temp(19989 downto 19980) := ADC(11 downto 2);
					when 1999 => temp(19999 downto 19990) := ADC(11 downto 2);
					when 2000 => temp(20009 downto 20000) := ADC(11 downto 2);
					when 2001 => temp(20019 downto 20010) := ADC(11 downto 2);
					when 2002 => temp(20029 downto 20020) := ADC(11 downto 2);
					when 2003 => temp(20039 downto 20030) := ADC(11 downto 2);
					when 2004 => temp(20049 downto 20040) := ADC(11 downto 2);
					when 2005 => temp(20059 downto 20050) := ADC(11 downto 2);
					when 2006 => temp(20069 downto 20060) := ADC(11 downto 2);
					when 2007 => temp(20079 downto 20070) := ADC(11 downto 2);
					when 2008 => temp(20089 downto 20080) := ADC(11 downto 2);
					when 2009 => temp(20099 downto 20090) := ADC(11 downto 2);
					when 2010 => temp(20109 downto 20100) := ADC(11 downto 2);
					when 2011 => temp(20119 downto 20110) := ADC(11 downto 2);
					when 2012 => temp(20129 downto 20120) := ADC(11 downto 2);
					when 2013 => temp(20139 downto 20130) := ADC(11 downto 2);
					when 2014 => temp(20149 downto 20140) := ADC(11 downto 2);
					when 2015 => temp(20159 downto 20150) := ADC(11 downto 2);
					when 2016 => temp(20169 downto 20160) := ADC(11 downto 2);
					when 2017 => temp(20179 downto 20170) := ADC(11 downto 2);
					when 2018 => temp(20189 downto 20180) := ADC(11 downto 2);
					when 2019 => temp(20199 downto 20190) := ADC(11 downto 2);
					when 2020 => temp(20209 downto 20200) := ADC(11 downto 2);
					when 2021 => temp(20219 downto 20210) := ADC(11 downto 2);
					when 2022 => temp(20229 downto 20220) := ADC(11 downto 2);
					when 2023 => temp(20239 downto 20230) := ADC(11 downto 2);
					when 2024 => temp(20249 downto 20240) := ADC(11 downto 2);
					when 2025 => temp(20259 downto 20250) := ADC(11 downto 2);
					when 2026 => temp(20269 downto 20260) := ADC(11 downto 2);
					when 2027 => temp(20279 downto 20270) := ADC(11 downto 2);
					when 2028 => temp(20289 downto 20280) := ADC(11 downto 2);
					when 2029 => temp(20299 downto 20290) := ADC(11 downto 2);
					when 2030 => temp(20309 downto 20300) := ADC(11 downto 2);
					when 2031 => temp(20319 downto 20310) := ADC(11 downto 2);
					when 2032 => temp(20329 downto 20320) := ADC(11 downto 2);
					when 2033 => temp(20339 downto 20330) := ADC(11 downto 2);
					when 2034 => temp(20349 downto 20340) := ADC(11 downto 2);
					when 2035 => temp(20359 downto 20350) := ADC(11 downto 2);
					when 2036 => temp(20369 downto 20360) := ADC(11 downto 2);
					when 2037 => temp(20379 downto 20370) := ADC(11 downto 2);
					when 2038 => temp(20389 downto 20380) := ADC(11 downto 2);
					when 2039 => temp(20399 downto 20390) := ADC(11 downto 2);
					when 2040 => temp(20409 downto 20400) := ADC(11 downto 2);
					when 2041 => temp(20419 downto 20410) := ADC(11 downto 2);
					when 2042 => temp(20429 downto 20420) := ADC(11 downto 2);
					when 2043 => temp(20439 downto 20430) := ADC(11 downto 2);
					when 2044 => temp(20449 downto 20440) := ADC(11 downto 2);
					when 2045 => temp(20459 downto 20450) := ADC(11 downto 2);
					when 2046 => temp(20469 downto 20460) := ADC(11 downto 2);
					when 2047 => temp(20479 downto 20470) := ADC(11 downto 2);
					when others => null;
					----------------------------------------
				end case;
					
--------------------------------------
-- state 4 increment             --
--------------------------------------
	when state_4 =>
					next_state <= state_2;
				--------------------------
				--  determine outputs   --
				--------------------------
				DONE			<= '1';
				ADC_CONVST	<= '1';
				ADC_WB		<= '1';
				ADC_WR		<= '1';
				ADC_RD		<= '1';
				ADC_CS		<= '0';
				ADC 			<= "ZZZZZZZZZZZZ";
				LEDG 			<= "00010000";
				timer_reset <= '1';
				setup_timer_reset <= '1';
				sample_counter_increment <= '1';
				sample_counter_reset <= '0';

--------------------------------------
-- state 5 done              		--
--------------------------------------
			when state_5 =>
				--------------------------
				-- determine next state --
				--------------------------
				if (CONTROL = '0')
				then
					next_state <= state_1;
				else
					next_state <= present_state;
				end if;
				--------------------------
				--  determine outputs   --
				--------------------------
				DONE			<= '1';
				ADC_CONVST	<= '1';
				ADC_WB		<= '1';
				ADC_WR		<= '1';
				ADC_RD		<= '1';
				ADC_CS		<= '0';
				ADC 			<= "ZZZZZZZZZZZZ";
				LEDG 			<= "00100000";
				timer_reset <= '1';
				setup_timer_reset <= '1';
				sample_counter_increment <= '0';
				sample_counter_reset <= '1';
--------------------------------------
--  unknown state returns to init   --
--------------------------------------
			when others =>
				next_state <= state_0;
		end case;

		samples <= temp;

	end process;
end ADC_sampler;