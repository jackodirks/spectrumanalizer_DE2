-- nios2VGA.vhd

-- Generated using ACDS version 13.0sp1 232 at 2014.01.20.12:59:07

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios2VGA is
	port (
		clk_clk                                  : in    std_logic                     := '0';             --                               clk.clk
		reset_reset_n                            : in    std_logic                     := '0';             --                             reset.reset_n
		red_led_pio_external_connection_export   : out   std_logic_vector(17 downto 0);                    --   red_led_pio_external_connection.export
		vga_controller_external_CLK              : out   std_logic;                                        --           vga_controller_external.CLK
		vga_controller_external_HS               : out   std_logic;                                        --                                  .HS
		vga_controller_external_VS               : out   std_logic;                                        --                                  .VS
		vga_controller_external_BLANK            : out   std_logic;                                        --                                  .BLANK
		vga_controller_external_SYNC             : out   std_logic;                                        --                                  .SYNC
		vga_controller_external_R                : out   std_logic_vector(9 downto 0);                     --                                  .R
		vga_controller_external_G                : out   std_logic_vector(9 downto 0);                     --                                  .G
		vga_controller_external_B                : out   std_logic_vector(9 downto 0);                     --                                  .B
		sram_external_interface_DQ               : inout std_logic_vector(15 downto 0) := (others => '0'); --           sram_external_interface.DQ
		sram_external_interface_ADDR             : out   std_logic_vector(17 downto 0);                    --                                  .ADDR
		sram_external_interface_LB_N             : out   std_logic;                                        --                                  .LB_N
		sram_external_interface_UB_N             : out   std_logic;                                        --                                  .UB_N
		sram_external_interface_CE_N             : out   std_logic;                                        --                                  .CE_N
		sram_external_interface_OE_N             : out   std_logic;                                        --                                  .OE_N
		sram_external_interface_WE_N             : out   std_logic;                                        --                                  .WE_N
		vga_clock_out_clk_clk                    : out   std_logic;                                        --                 vga_clock_out_clk.clk
		green_led_pio_external_connection_export : out   std_logic_vector(8 downto 0);                     -- green_led_pio_external_connection.export
		sdram_clock_clk                          : out   std_logic;                                        --                       sdram_clock.clk
		nios_cntrl_in_export                     : in    std_logic_vector(7 downto 0)  := (others => '0'); --                     nios_cntrl_in.export
		nios_cntrl_out_export                    : out   std_logic_vector(7 downto 0);                     --                    nios_cntrl_out.export
		fft_in_0_export                          : in    std_logic_vector(31 downto 0) := (others => '0'); --                          fft_in_0.export
		fft_in_1_export                          : in    std_logic_vector(31 downto 0) := (others => '0'); --                          fft_in_1.export
		fft_in_2_export                          : in    std_logic_vector(31 downto 0) := (others => '0'); --                          fft_in_2.export
		fft_in_3_export                          : in    std_logic_vector(31 downto 0) := (others => '0'); --                          fft_in_3.export
		rotary_in_export                         : in    std_logic_vector(7 downto 0)  := (others => '0')  --                         rotary_in.export
	);
end entity nios2VGA;

architecture rtl of nios2VGA is
	component nios2VGA_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(19 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios2VGA_cpu;

	component nios2VGA_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios2VGA_jtag_uart;

	component nios2VGA_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios2VGA_sys_clk_timer;

	component nios2VGA_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios2VGA_sysid;

	component nios2VGA_red_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component nios2VGA_red_led_pio;

	component nios2VGA_external_clocks is
		port (
			CLOCK_50    : in  std_logic := 'X'; -- clk
			reset       : in  std_logic := 'X'; -- reset
			sys_clk     : out std_logic;        -- clk
			sys_reset_n : out std_logic;        -- reset_n
			SDRAM_CLK   : out std_logic;        -- clk
			VGA_CLK     : out std_logic         -- clk
		);
	end component nios2VGA_external_clocks;

	component nios2VGA_VGA_Dual_Clock_FIFO is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component nios2VGA_VGA_Dual_Clock_FIFO;

	component nios2VGA_Alpha_Blending is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			foreground_data          : in  std_logic_vector(39 downto 0) := (others => 'X'); -- data
			foreground_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			foreground_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			foreground_valid         : in  std_logic                     := 'X';             -- valid
			foreground_ready         : out std_logic;                                        -- ready
			background_data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			background_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			background_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			background_valid         : in  std_logic                     := 'X';             -- valid
			background_ready         : out std_logic;                                        -- ready
			output_ready             : in  std_logic                     := 'X';             -- ready
			output_data              : out std_logic_vector(29 downto 0);                    -- data
			output_startofpacket     : out std_logic;                                        -- startofpacket
			output_endofpacket       : out std_logic;                                        -- endofpacket
			output_valid             : out std_logic                                         -- valid
		);
	end component nios2VGA_Alpha_Blending;

	component nios2VGA_VGA_Controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(9 downto 0);                     -- export
			VGA_G         : out std_logic_vector(9 downto 0);                     -- export
			VGA_B         : out std_logic_vector(9 downto 0)                      -- export
		);
	end component nios2VGA_VGA_Controller;

	component nios2VGA_VGA_Character_buffer is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			ctrl_address         : in  std_logic                     := 'X';             -- address
			ctrl_byteenable      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ctrl_chipselect      : in  std_logic                     := 'X';             -- chipselect
			ctrl_read            : in  std_logic                     := 'X';             -- read
			ctrl_write           : in  std_logic                     := 'X';             -- write
			ctrl_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ctrl_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			buf_byteenable       : in  std_logic                     := 'X';             -- byteenable
			buf_chipselect       : in  std_logic                     := 'X';             -- chipselect
			buf_read             : in  std_logic                     := 'X';             -- read
			buf_write            : in  std_logic                     := 'X';             -- write
			buf_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			buf_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			buf_waitrequest      : out std_logic;                                        -- waitrequest
			buf_address          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(39 downto 0)                     -- data
		);
	end component nios2VGA_VGA_Character_buffer;

	component nios2VGA_VGA_Scaler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component nios2VGA_VGA_Scaler;

	component nios2VGA_VGA_pixel_RGB_Resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component nios2VGA_VGA_pixel_RGB_Resampler;

	component nios2VGA_VGA_Pixel_Buffer is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component nios2VGA_VGA_Pixel_Buffer;

	component nios2VGA_SRAM is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(17 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(17 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component nios2VGA_SRAM;

	component nios2VGA_green_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component nios2VGA_green_led_pio;

	component nios2VGA_control_in is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component nios2VGA_control_in;

	component nios2VGA_control_out is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios2VGA_control_out;

	component nios2VGA_FFT_in_0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component nios2VGA_FFT_in_0;

	component nios2VGA_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios2VGA_addr_router;

	component nios2VGA_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(90 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2VGA_addr_router_001;

	component nios2VGA_addr_router_002 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios2VGA_addr_router_002;

	component nios2VGA_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios2VGA_id_router;

	component nios2VGA_id_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(90 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2VGA_id_router_001;

	component nios2VGA_id_router_002 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios2VGA_id_router_002;

	component nios2VGA_id_router_007 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(81 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios2VGA_id_router_007;

	component nios2VGA_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(108 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(108 downto 0);                    -- data
			src1_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component nios2VGA_cmd_xbar_demux;

	component nios2VGA_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(90 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios2VGA_cmd_xbar_demux_001;

	component nios2VGA_cmd_xbar_demux_002 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			sink_ready          : out std_logic;                                         -- ready
			sink_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready          : in  std_logic                      := 'X';             -- ready
			src0_valid          : out std_logic;                                         -- valid
			src0_data           : out std_logic_vector(108 downto 0);                    -- data
			src0_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src0_startofpacket  : out std_logic;                                         -- startofpacket
			src0_endofpacket    : out std_logic;                                         -- endofpacket
			src1_ready          : in  std_logic                      := 'X';             -- ready
			src1_valid          : out std_logic;                                         -- valid
			src1_data           : out std_logic_vector(108 downto 0);                    -- data
			src1_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src1_startofpacket  : out std_logic;                                         -- startofpacket
			src1_endofpacket    : out std_logic;                                         -- endofpacket
			src2_ready          : in  std_logic                      := 'X';             -- ready
			src2_valid          : out std_logic;                                         -- valid
			src2_data           : out std_logic_vector(108 downto 0);                    -- data
			src2_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src2_startofpacket  : out std_logic;                                         -- startofpacket
			src2_endofpacket    : out std_logic;                                         -- endofpacket
			src3_ready          : in  std_logic                      := 'X';             -- ready
			src3_valid          : out std_logic;                                         -- valid
			src3_data           : out std_logic_vector(108 downto 0);                    -- data
			src3_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src3_startofpacket  : out std_logic;                                         -- startofpacket
			src3_endofpacket    : out std_logic;                                         -- endofpacket
			src4_ready          : in  std_logic                      := 'X';             -- ready
			src4_valid          : out std_logic;                                         -- valid
			src4_data           : out std_logic_vector(108 downto 0);                    -- data
			src4_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src4_startofpacket  : out std_logic;                                         -- startofpacket
			src4_endofpacket    : out std_logic;                                         -- endofpacket
			src5_ready          : in  std_logic                      := 'X';             -- ready
			src5_valid          : out std_logic;                                         -- valid
			src5_data           : out std_logic_vector(108 downto 0);                    -- data
			src5_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src5_startofpacket  : out std_logic;                                         -- startofpacket
			src5_endofpacket    : out std_logic;                                         -- endofpacket
			src6_ready          : in  std_logic                      := 'X';             -- ready
			src6_valid          : out std_logic;                                         -- valid
			src6_data           : out std_logic_vector(108 downto 0);                    -- data
			src6_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src6_startofpacket  : out std_logic;                                         -- startofpacket
			src6_endofpacket    : out std_logic;                                         -- endofpacket
			src7_ready          : in  std_logic                      := 'X';             -- ready
			src7_valid          : out std_logic;                                         -- valid
			src7_data           : out std_logic_vector(108 downto 0);                    -- data
			src7_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src7_startofpacket  : out std_logic;                                         -- startofpacket
			src7_endofpacket    : out std_logic;                                         -- endofpacket
			src8_ready          : in  std_logic                      := 'X';             -- ready
			src8_valid          : out std_logic;                                         -- valid
			src8_data           : out std_logic_vector(108 downto 0);                    -- data
			src8_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src8_startofpacket  : out std_logic;                                         -- startofpacket
			src8_endofpacket    : out std_logic;                                         -- endofpacket
			src9_ready          : in  std_logic                      := 'X';             -- ready
			src9_valid          : out std_logic;                                         -- valid
			src9_data           : out std_logic_vector(108 downto 0);                    -- data
			src9_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src9_startofpacket  : out std_logic;                                         -- startofpacket
			src9_endofpacket    : out std_logic;                                         -- endofpacket
			src10_ready         : in  std_logic                      := 'X';             -- ready
			src10_valid         : out std_logic;                                         -- valid
			src10_data          : out std_logic_vector(108 downto 0);                    -- data
			src10_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src10_startofpacket : out std_logic;                                         -- startofpacket
			src10_endofpacket   : out std_logic;                                         -- endofpacket
			src11_ready         : in  std_logic                      := 'X';             -- ready
			src11_valid         : out std_logic;                                         -- valid
			src11_data          : out std_logic_vector(108 downto 0);                    -- data
			src11_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src11_startofpacket : out std_logic;                                         -- startofpacket
			src11_endofpacket   : out std_logic;                                         -- endofpacket
			src12_ready         : in  std_logic                      := 'X';             -- ready
			src12_valid         : out std_logic;                                         -- valid
			src12_data          : out std_logic_vector(108 downto 0);                    -- data
			src12_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src12_startofpacket : out std_logic;                                         -- startofpacket
			src12_endofpacket   : out std_logic;                                         -- endofpacket
			src13_ready         : in  std_logic                      := 'X';             -- ready
			src13_valid         : out std_logic;                                         -- valid
			src13_data          : out std_logic_vector(108 downto 0);                    -- data
			src13_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src13_startofpacket : out std_logic;                                         -- startofpacket
			src13_endofpacket   : out std_logic;                                         -- endofpacket
			src14_ready         : in  std_logic                      := 'X';             -- ready
			src14_valid         : out std_logic;                                         -- valid
			src14_data          : out std_logic_vector(108 downto 0);                    -- data
			src14_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src14_startofpacket : out std_logic;                                         -- startofpacket
			src14_endofpacket   : out std_logic;                                         -- endofpacket
			src15_ready         : in  std_logic                      := 'X';             -- ready
			src15_valid         : out std_logic;                                         -- valid
			src15_data          : out std_logic_vector(108 downto 0);                    -- data
			src15_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src15_startofpacket : out std_logic;                                         -- startofpacket
			src15_endofpacket   : out std_logic;                                         -- endofpacket
			src16_ready         : in  std_logic                      := 'X';             -- ready
			src16_valid         : out std_logic;                                         -- valid
			src16_data          : out std_logic_vector(108 downto 0);                    -- data
			src16_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src16_startofpacket : out std_logic;                                         -- startofpacket
			src16_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component nios2VGA_cmd_xbar_demux_002;

	component nios2VGA_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(108 downto 0);                    -- data
			src_channel         : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component nios2VGA_cmd_xbar_mux;

	component nios2VGA_cmd_xbar_mux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(90 downto 0);                    -- data
			src_channel         : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios2VGA_cmd_xbar_mux_001;

	component nios2VGA_rsp_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(90 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(90 downto 0);                    -- data
			src1_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(90 downto 0);                    -- data
			src2_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios2VGA_rsp_xbar_demux_001;

	component nios2VGA_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(108 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component nios2VGA_rsp_xbar_demux_002;

	component nios2VGA_rsp_xbar_demux_007 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(81 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios2VGA_rsp_xbar_demux_007;

	component nios2VGA_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(108 downto 0);                    -- data
			src_channel         : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component nios2VGA_rsp_xbar_mux;

	component nios2VGA_rsp_xbar_mux_002 is
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			src_ready            : in  std_logic                      := 'X';             -- ready
			src_valid            : out std_logic;                                         -- valid
			src_data             : out std_logic_vector(108 downto 0);                    -- data
			src_channel          : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket    : out std_logic;                                         -- startofpacket
			src_endofpacket      : out std_logic;                                         -- endofpacket
			sink0_ready          : out std_logic;                                         -- ready
			sink0_valid          : in  std_logic                      := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                         -- ready
			sink1_valid          : in  std_logic                      := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                         -- ready
			sink2_valid          : in  std_logic                      := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                         -- ready
			sink3_valid          : in  std_logic                      := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                         -- ready
			sink4_valid          : in  std_logic                      := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                         -- ready
			sink5_valid          : in  std_logic                      := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                         -- ready
			sink6_valid          : in  std_logic                      := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                         -- ready
			sink7_valid          : in  std_logic                      := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                         -- ready
			sink8_valid          : in  std_logic                      := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                         -- ready
			sink9_valid          : in  std_logic                      := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                         -- ready
			sink10_valid         : in  std_logic                      := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                         -- ready
			sink11_valid         : in  std_logic                      := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                         -- ready
			sink12_valid         : in  std_logic                      := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                         -- ready
			sink13_valid         : in  std_logic                      := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink14_ready         : out std_logic;                                         -- ready
			sink14_valid         : in  std_logic                      := 'X';             -- valid
			sink14_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink14_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink14_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink14_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink15_ready         : out std_logic;                                         -- ready
			sink15_valid         : in  std_logic                      := 'X';             -- valid
			sink15_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink15_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink15_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink15_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink16_ready         : out std_logic;                                         -- ready
			sink16_valid         : in  std_logic                      := 'X';             -- valid
			sink16_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink16_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink16_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink16_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component nios2VGA_rsp_xbar_mux_002;

	component nios2VGA_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios2VGA_irq_mapper;

	component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(109 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(109 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(33 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(91 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(91 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(82 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(9 downto 0);                     -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(108 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(109 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(109 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(90 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(91 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(91 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent;

	component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(0 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(7 downto 0);                     -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(81 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(82 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(9 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent;

	component nios2vga_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(90 downto 0);                     -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component nios2vga_width_adapter;

	component nios2vga_width_adapter_002 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(81 downto 0);                     -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component nios2vga_width_adapter_002;

	component nios2vga_width_adapter_003 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(90 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(108 downto 0);                    -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component nios2vga_width_adapter_003;

	component nios2vga_width_adapter_005 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(81 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(108 downto 0);                    -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component nios2vga_width_adapter_005;

	component nios2vga_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios2vga_cpu_instruction_master_translator;

	component nios2vga_vga_pixel_buffer_avalon_pixel_dma_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(15 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios2vga_vga_pixel_buffer_avalon_pixel_dma_master_translator;

	component nios2vga_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios2vga_cpu_data_master_translator;

	component nios2vga_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(90 downto 0);                    -- data
			source0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component nios2vga_burst_adapter;

	component nios2vga_burst_adapter_001 is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(81 downto 0);                    -- data
			source0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component nios2vga_burst_adapter_001;

	component nios2vga_crosser is
		generic (
			DATA_WIDTH          : integer := 8;
			BITS_PER_SYMBOL     : integer := 8;
			USE_PACKETS         : integer := 0;
			USE_CHANNEL         : integer := 0;
			CHANNEL_WIDTH       : integer := 1;
			USE_ERROR           : integer := 0;
			ERROR_WIDTH         : integer := 1;
			VALID_SYNC_DEPTH    : integer := 2;
			READY_SYNC_DEPTH    : integer := 2;
			USE_OUTPUT_PIPELINE : integer := 1
		);
		port (
			in_clk            : in  std_logic                      := 'X';             -- clk
			in_reset          : in  std_logic                      := 'X';             -- reset
			out_clk           : in  std_logic                      := 'X';             -- clk
			out_reset         : in  std_logic                      := 'X';             -- reset
			in_ready          : out std_logic;                                         -- ready
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_valid         : out std_logic;                                         -- valid
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_channel       : out std_logic_vector(16 downto 0);                     -- channel
			out_data          : out std_logic_vector(108 downto 0);                    -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_empty         : out std_logic;                                         -- empty
			out_error         : out std_logic                                          -- error
		);
	end component nios2vga_crosser;

	component nios2vga_crosser_004 is
		generic (
			DATA_WIDTH          : integer := 8;
			BITS_PER_SYMBOL     : integer := 8;
			USE_PACKETS         : integer := 0;
			USE_CHANNEL         : integer := 0;
			CHANNEL_WIDTH       : integer := 1;
			USE_ERROR           : integer := 0;
			ERROR_WIDTH         : integer := 1;
			VALID_SYNC_DEPTH    : integer := 2;
			READY_SYNC_DEPTH    : integer := 2;
			USE_OUTPUT_PIPELINE : integer := 1
		);
		port (
			in_clk            : in  std_logic                     := 'X';             -- clk
			in_reset          : in  std_logic                     := 'X';             -- reset
			out_clk           : in  std_logic                     := 'X';             -- clk
			out_reset         : in  std_logic                     := 'X';             -- reset
			in_ready          : out std_logic;                                        -- ready
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_channel        : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			in_data           : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_valid         : out std_logic;                                        -- valid
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			out_channel       : out std_logic_vector(16 downto 0);                    -- channel
			out_data          : out std_logic_vector(90 downto 0);                    -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_empty         : out std_logic;                                        -- empty
			out_error         : out std_logic                                         -- error
		);
	end component nios2vga_crosser_004;

	component nios2vga_crosser_006 is
		generic (
			DATA_WIDTH          : integer := 8;
			BITS_PER_SYMBOL     : integer := 8;
			USE_PACKETS         : integer := 0;
			USE_CHANNEL         : integer := 0;
			CHANNEL_WIDTH       : integer := 1;
			USE_ERROR           : integer := 0;
			ERROR_WIDTH         : integer := 1;
			VALID_SYNC_DEPTH    : integer := 2;
			READY_SYNC_DEPTH    : integer := 2;
			USE_OUTPUT_PIPELINE : integer := 1
		);
		port (
			in_clk            : in  std_logic                     := 'X';             -- clk
			in_reset          : in  std_logic                     := 'X';             -- reset
			out_clk           : in  std_logic                     := 'X';             -- clk
			out_reset         : in  std_logic                     := 'X';             -- reset
			in_ready          : out std_logic;                                        -- ready
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_channel        : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			in_data           : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_valid         : out std_logic;                                        -- valid
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			out_channel       : out std_logic_vector(16 downto 0);                    -- channel
			out_data          : out std_logic_vector(81 downto 0);                    -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_empty         : out std_logic;                                        -- empty
			out_error         : out std_logic                                         -- error
		);
	end component nios2vga_crosser_006;

	component nios2vga_cpu_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_cpu_jtag_debug_module_translator;

	component nios2vga_sram_avalon_sram_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(17 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_sram_avalon_sram_slave_translator;

	component nios2vga_jtag_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_jtag_uart_avalon_jtag_slave_translator;

	component nios2vga_sys_clk_timer_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_sys_clk_timer_s1_translator;

	component nios2vga_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_sysid_control_slave_translator;

	component nios2vga_red_led_pio_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_red_led_pio_s1_translator;

	component nios2vga_vga_character_buffer_avalon_char_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_vga_character_buffer_avalon_char_control_slave_translator;

	component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(7 downto 0);                     -- readdata
			uav_writedata            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(12 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator;

	component nios2vga_vga_pixel_buffer_avalon_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_vga_pixel_buffer_avalon_control_slave_translator;

	component nios2vga_control_in_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios2vga_control_in_s1_translator;

	component nios2vga_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component nios2vga_rst_controller;

	component nios2vga_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component nios2vga_rst_controller_001;

	component nios2vga_cpu_instruction_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(108 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component nios2vga_cpu_instruction_master_translator_avalon_universal_master_0_agent;

	component nios2vga_vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(90 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component nios2vga_vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent;

	signal external_clocks_vga_clk_clk                                                                                         : std_logic;                      -- external_clocks:VGA_CLK -> [vga_clock_out_clk_clk, VGA_Controller:clk, VGA_Dual_Clock_FIFO:clk_stream_out, rst_controller_003:clk]
	signal external_clocks_sys_clk_clk                                                                                         : std_logic;                      -- external_clocks:sys_clk -> [Alpha_Blending:clk, SRAM:clk, SRAM_avalon_sram_slave_translator:clk, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Character_buffer:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Character_buffer_avalon_char_control_slave_translator:clk, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:clk, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Dual_Clock_FIFO:clk_stream_in, VGA_Pixel_Buffer:clk, VGA_Pixel_Buffer_avalon_control_slave_translator:clk, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:clk, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, VGA_Scaler:clk, VGA_pixel_RGB_Resampler:clk, addr_router_001:clk, burst_adapter:clk, burst_adapter_001:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux_001:clk, crosser:out_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, crosser_004:out_clk, crosser_005:out_clk, crosser_006:out_clk, crosser_007:in_clk, crosser_008:in_clk, crosser_009:in_clk, id_router_001:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rst_controller_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk]
	signal vga_character_buffer_avalon_char_source_endofpacket                                                                 : std_logic;                      -- VGA_Character_buffer:stream_endofpacket -> Alpha_Blending:foreground_endofpacket
	signal vga_character_buffer_avalon_char_source_valid                                                                       : std_logic;                      -- VGA_Character_buffer:stream_valid -> Alpha_Blending:foreground_valid
	signal vga_character_buffer_avalon_char_source_startofpacket                                                               : std_logic;                      -- VGA_Character_buffer:stream_startofpacket -> Alpha_Blending:foreground_startofpacket
	signal vga_character_buffer_avalon_char_source_data                                                                        : std_logic_vector(39 downto 0);  -- VGA_Character_buffer:stream_data -> Alpha_Blending:foreground_data
	signal vga_character_buffer_avalon_char_source_ready                                                                       : std_logic;                      -- Alpha_Blending:foreground_ready -> VGA_Character_buffer:stream_ready
	signal alpha_blending_avalon_blended_source_endofpacket                                                                    : std_logic;                      -- Alpha_Blending:output_endofpacket -> VGA_Dual_Clock_FIFO:stream_in_endofpacket
	signal alpha_blending_avalon_blended_source_valid                                                                          : std_logic;                      -- Alpha_Blending:output_valid -> VGA_Dual_Clock_FIFO:stream_in_valid
	signal alpha_blending_avalon_blended_source_startofpacket                                                                  : std_logic;                      -- Alpha_Blending:output_startofpacket -> VGA_Dual_Clock_FIFO:stream_in_startofpacket
	signal alpha_blending_avalon_blended_source_data                                                                           : std_logic_vector(29 downto 0);  -- Alpha_Blending:output_data -> VGA_Dual_Clock_FIFO:stream_in_data
	signal alpha_blending_avalon_blended_source_ready                                                                          : std_logic;                      -- VGA_Dual_Clock_FIFO:stream_in_ready -> Alpha_Blending:output_ready
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket                                                             : std_logic;                      -- VGA_Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_valid                                                                   : std_logic;                      -- VGA_Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket                                                           : std_logic;                      -- VGA_Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_data                                                                    : std_logic_vector(29 downto 0);  -- VGA_Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_ready                                                                   : std_logic;                      -- VGA_Controller:ready -> VGA_Dual_Clock_FIFO:stream_out_ready
	signal vga_scaler_avalon_scaler_source_endofpacket                                                                         : std_logic;                      -- VGA_Scaler:stream_out_endofpacket -> Alpha_Blending:background_endofpacket
	signal vga_scaler_avalon_scaler_source_valid                                                                               : std_logic;                      -- VGA_Scaler:stream_out_valid -> Alpha_Blending:background_valid
	signal vga_scaler_avalon_scaler_source_startofpacket                                                                       : std_logic;                      -- VGA_Scaler:stream_out_startofpacket -> Alpha_Blending:background_startofpacket
	signal vga_scaler_avalon_scaler_source_data                                                                                : std_logic_vector(29 downto 0);  -- VGA_Scaler:stream_out_data -> Alpha_Blending:background_data
	signal vga_scaler_avalon_scaler_source_ready                                                                               : std_logic;                      -- Alpha_Blending:background_ready -> VGA_Scaler:stream_out_ready
	signal vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket                                                               : std_logic;                      -- VGA_pixel_RGB_Resampler:stream_out_endofpacket -> VGA_Scaler:stream_in_endofpacket
	signal vga_pixel_rgb_resampler_avalon_rgb_source_valid                                                                     : std_logic;                      -- VGA_pixel_RGB_Resampler:stream_out_valid -> VGA_Scaler:stream_in_valid
	signal vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket                                                             : std_logic;                      -- VGA_pixel_RGB_Resampler:stream_out_startofpacket -> VGA_Scaler:stream_in_startofpacket
	signal vga_pixel_rgb_resampler_avalon_rgb_source_data                                                                      : std_logic_vector(29 downto 0);  -- VGA_pixel_RGB_Resampler:stream_out_data -> VGA_Scaler:stream_in_data
	signal vga_pixel_rgb_resampler_avalon_rgb_source_ready                                                                     : std_logic;                      -- VGA_Scaler:stream_in_ready -> VGA_pixel_RGB_Resampler:stream_out_ready
	signal vga_pixel_buffer_avalon_pixel_source_endofpacket                                                                    : std_logic;                      -- VGA_Pixel_Buffer:stream_endofpacket -> VGA_pixel_RGB_Resampler:stream_in_endofpacket
	signal vga_pixel_buffer_avalon_pixel_source_valid                                                                          : std_logic;                      -- VGA_Pixel_Buffer:stream_valid -> VGA_pixel_RGB_Resampler:stream_in_valid
	signal vga_pixel_buffer_avalon_pixel_source_startofpacket                                                                  : std_logic;                      -- VGA_Pixel_Buffer:stream_startofpacket -> VGA_pixel_RGB_Resampler:stream_in_startofpacket
	signal vga_pixel_buffer_avalon_pixel_source_data                                                                           : std_logic_vector(15 downto 0);  -- VGA_Pixel_Buffer:stream_data -> VGA_pixel_RGB_Resampler:stream_in_data
	signal vga_pixel_buffer_avalon_pixel_source_ready                                                                          : std_logic;                      -- VGA_pixel_RGB_Resampler:stream_in_ready -> VGA_Pixel_Buffer:stream_ready
	signal cpu_instruction_master_waitrequest                                                                                  : std_logic;                      -- cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                                                                      : std_logic_vector(19 downto 0);  -- cpu:i_address -> cpu_instruction_master_translator:av_address
	signal cpu_instruction_master_read                                                                                         : std_logic;                      -- cpu:i_read -> cpu_instruction_master_translator:av_read
	signal cpu_instruction_master_readdata                                                                                     : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	signal vga_pixel_buffer_avalon_pixel_dma_master_waitrequest                                                                : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_waitrequest -> VGA_Pixel_Buffer:master_waitrequest
	signal vga_pixel_buffer_avalon_pixel_dma_master_address                                                                    : std_logic_vector(31 downto 0);  -- VGA_Pixel_Buffer:master_address -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_address
	signal vga_pixel_buffer_avalon_pixel_dma_master_lock                                                                       : std_logic;                      -- VGA_Pixel_Buffer:master_arbiterlock -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_lock
	signal vga_pixel_buffer_avalon_pixel_dma_master_read                                                                       : std_logic;                      -- VGA_Pixel_Buffer:master_read -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_read
	signal vga_pixel_buffer_avalon_pixel_dma_master_readdata                                                                   : std_logic_vector(15 downto 0);  -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_readdata -> VGA_Pixel_Buffer:master_readdata
	signal vga_pixel_buffer_avalon_pixel_dma_master_readdatavalid                                                              : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_readdatavalid -> VGA_Pixel_Buffer:master_readdatavalid
	signal cpu_data_master_waitrequest                                                                                         : std_logic;                      -- cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_writedata                                                                                           : std_logic_vector(31 downto 0);  -- cpu:d_writedata -> cpu_data_master_translator:av_writedata
	signal cpu_data_master_address                                                                                             : std_logic_vector(19 downto 0);  -- cpu:d_address -> cpu_data_master_translator:av_address
	signal cpu_data_master_write                                                                                               : std_logic;                      -- cpu:d_write -> cpu_data_master_translator:av_write
	signal cpu_data_master_read                                                                                                : std_logic;                      -- cpu:d_read -> cpu_data_master_translator:av_read
	signal cpu_data_master_readdata                                                                                            : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:av_readdata -> cpu:d_readdata
	signal cpu_data_master_debugaccess                                                                                         : std_logic;                      -- cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	signal cpu_data_master_byteenable                                                                                          : std_logic_vector(3 downto 0);   -- cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                                    : std_logic;                      -- cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                                      : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_address                                                        : std_logic_vector(8 downto 0);   -- cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_write                                                          : std_logic;                      -- cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_read                                                           : std_logic;                      -- cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                                       : std_logic_vector(31 downto 0);  -- cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                                    : std_logic;                      -- cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                                     : std_logic_vector(3 downto 0);   -- cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(15 downto 0);  -- SRAM_avalon_sram_slave_translator:av_writedata -> SRAM:writedata
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(17 downto 0);  -- SRAM_avalon_sram_slave_translator:av_address -> SRAM:address
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- SRAM_avalon_sram_slave_translator:av_write -> SRAM:write
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_read                                                          : std_logic;                      -- SRAM_avalon_sram_slave_translator:av_read -> SRAM:read
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(15 downto 0);  -- SRAM:readdata -> SRAM_avalon_sram_slave_translator:av_readdata
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid                                                 : std_logic;                      -- SRAM:readdatavalid -> SRAM_avalon_sram_slave_translator:av_readdatavalid
	signal sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable                                                    : std_logic_vector(1 downto 0);   -- SRAM_avalon_sram_slave_translator:av_byteenable -> SRAM:byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                                              : std_logic;                      -- jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(0 downto 0);   -- jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                                    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                                     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata                                                           : std_logic_vector(15 downto 0);  -- sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_address                                                             : std_logic_vector(2 downto 0);   -- sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect                                                          : std_logic;                      -- sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_write                                                               : std_logic;                      -- sys_clk_timer_s1_translator:av_write -> sys_clk_timer_s1_translator_avalon_anti_slave_0_write:in
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata                                                            : std_logic_vector(15 downto 0);  -- sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                                          : std_logic_vector(0 downto 0);   -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                                         : std_logic_vector(31 downto 0);  -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal red_led_pio_s1_translator_avalon_anti_slave_0_writedata                                                             : std_logic_vector(31 downto 0);  -- red_led_pio_s1_translator:av_writedata -> red_led_pio:writedata
	signal red_led_pio_s1_translator_avalon_anti_slave_0_address                                                               : std_logic_vector(1 downto 0);   -- red_led_pio_s1_translator:av_address -> red_led_pio:address
	signal red_led_pio_s1_translator_avalon_anti_slave_0_chipselect                                                            : std_logic;                      -- red_led_pio_s1_translator:av_chipselect -> red_led_pio:chipselect
	signal red_led_pio_s1_translator_avalon_anti_slave_0_write                                                                 : std_logic;                      -- red_led_pio_s1_translator:av_write -> red_led_pio_s1_translator_avalon_anti_slave_0_write:in
	signal red_led_pio_s1_translator_avalon_anti_slave_0_readdata                                                              : std_logic_vector(31 downto 0);  -- red_led_pio:readdata -> red_led_pio_s1_translator:av_readdata
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- VGA_Character_buffer_avalon_char_control_slave_translator:av_writedata -> VGA_Character_buffer:ctrl_writedata
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(0 downto 0);   -- VGA_Character_buffer_avalon_char_control_slave_translator:av_address -> VGA_Character_buffer:ctrl_address
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect                            : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator:av_chipselect -> VGA_Character_buffer:ctrl_chipselect
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator:av_write -> VGA_Character_buffer:ctrl_write
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator:av_read -> VGA_Character_buffer:ctrl_read
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- VGA_Character_buffer:ctrl_readdata -> VGA_Character_buffer_avalon_char_control_slave_translator:av_readdata
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- VGA_Character_buffer_avalon_char_control_slave_translator:av_byteenable -> VGA_Character_buffer:ctrl_byteenable
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest                            : std_logic;                      -- VGA_Character_buffer:buf_waitrequest -> VGA_Character_buffer_avalon_char_buffer_slave_translator:av_waitrequest
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(7 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator:av_writedata -> VGA_Character_buffer:buf_writedata
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address                                : std_logic_vector(12 downto 0);  -- VGA_Character_buffer_avalon_char_buffer_slave_translator:av_address -> VGA_Character_buffer:buf_address
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect                             : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator:av_chipselect -> VGA_Character_buffer:buf_chipselect
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write                                  : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator:av_write -> VGA_Character_buffer:buf_write
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read                                   : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator:av_read -> VGA_Character_buffer:buf_read
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(7 downto 0);   -- VGA_Character_buffer:buf_readdata -> VGA_Character_buffer_avalon_char_buffer_slave_translator:av_readdata
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable                             : std_logic_vector(0 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator:av_byteenable -> VGA_Character_buffer:buf_byteenable
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_writedata                                      : std_logic_vector(31 downto 0);  -- VGA_Pixel_Buffer_avalon_control_slave_translator:av_writedata -> VGA_Pixel_Buffer:slave_writedata
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_address                                        : std_logic_vector(1 downto 0);   -- VGA_Pixel_Buffer_avalon_control_slave_translator:av_address -> VGA_Pixel_Buffer:slave_address
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_write                                          : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator:av_write -> VGA_Pixel_Buffer:slave_write
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_read                                           : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator:av_read -> VGA_Pixel_Buffer:slave_read
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0);  -- VGA_Pixel_Buffer:slave_readdata -> VGA_Pixel_Buffer_avalon_control_slave_translator:av_readdata
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_byteenable                                     : std_logic_vector(3 downto 0);   -- VGA_Pixel_Buffer_avalon_control_slave_translator:av_byteenable -> VGA_Pixel_Buffer:slave_byteenable
	signal green_led_pio_s1_translator_avalon_anti_slave_0_writedata                                                           : std_logic_vector(31 downto 0);  -- green_led_pio_s1_translator:av_writedata -> green_led_pio:writedata
	signal green_led_pio_s1_translator_avalon_anti_slave_0_address                                                             : std_logic_vector(1 downto 0);   -- green_led_pio_s1_translator:av_address -> green_led_pio:address
	signal green_led_pio_s1_translator_avalon_anti_slave_0_chipselect                                                          : std_logic;                      -- green_led_pio_s1_translator:av_chipselect -> green_led_pio:chipselect
	signal green_led_pio_s1_translator_avalon_anti_slave_0_write                                                               : std_logic;                      -- green_led_pio_s1_translator:av_write -> green_led_pio_s1_translator_avalon_anti_slave_0_write:in
	signal green_led_pio_s1_translator_avalon_anti_slave_0_readdata                                                            : std_logic_vector(31 downto 0);  -- green_led_pio:readdata -> green_led_pio_s1_translator:av_readdata
	signal control_in_s1_translator_avalon_anti_slave_0_address                                                                : std_logic_vector(1 downto 0);   -- control_in_s1_translator:av_address -> control_in:address
	signal control_in_s1_translator_avalon_anti_slave_0_readdata                                                               : std_logic_vector(31 downto 0);  -- control_in:readdata -> control_in_s1_translator:av_readdata
	signal control_out_s1_translator_avalon_anti_slave_0_writedata                                                             : std_logic_vector(31 downto 0);  -- control_out_s1_translator:av_writedata -> control_out:writedata
	signal control_out_s1_translator_avalon_anti_slave_0_address                                                               : std_logic_vector(1 downto 0);   -- control_out_s1_translator:av_address -> control_out:address
	signal control_out_s1_translator_avalon_anti_slave_0_chipselect                                                            : std_logic;                      -- control_out_s1_translator:av_chipselect -> control_out:chipselect
	signal control_out_s1_translator_avalon_anti_slave_0_write                                                                 : std_logic;                      -- control_out_s1_translator:av_write -> control_out_s1_translator_avalon_anti_slave_0_write:in
	signal control_out_s1_translator_avalon_anti_slave_0_readdata                                                              : std_logic_vector(31 downto 0);  -- control_out:readdata -> control_out_s1_translator:av_readdata
	signal fft_in_0_s1_translator_avalon_anti_slave_0_address                                                                  : std_logic_vector(1 downto 0);   -- FFT_in_0_s1_translator:av_address -> FFT_in_0:address
	signal fft_in_0_s1_translator_avalon_anti_slave_0_readdata                                                                 : std_logic_vector(31 downto 0);  -- FFT_in_0:readdata -> FFT_in_0_s1_translator:av_readdata
	signal fft_in_1_s1_translator_avalon_anti_slave_0_address                                                                  : std_logic_vector(1 downto 0);   -- FFT_in_1_s1_translator:av_address -> FFT_in_1:address
	signal fft_in_1_s1_translator_avalon_anti_slave_0_readdata                                                                 : std_logic_vector(31 downto 0);  -- FFT_in_1:readdata -> FFT_in_1_s1_translator:av_readdata
	signal fft_in_2_s1_translator_avalon_anti_slave_0_address                                                                  : std_logic_vector(1 downto 0);   -- FFT_in_2_s1_translator:av_address -> FFT_in_2:address
	signal fft_in_2_s1_translator_avalon_anti_slave_0_readdata                                                                 : std_logic_vector(31 downto 0);  -- FFT_in_2:readdata -> FFT_in_2_s1_translator:av_readdata
	signal fft_in_3_s1_translator_avalon_anti_slave_0_address                                                                  : std_logic_vector(1 downto 0);   -- FFT_in_3_s1_translator:av_address -> FFT_in_3:address
	signal fft_in_3_s1_translator_avalon_anti_slave_0_readdata                                                                 : std_logic_vector(31 downto 0);  -- FFT_in_3:readdata -> FFT_in_3_s1_translator:av_readdata
	signal rotary_in_s1_translator_avalon_anti_slave_0_address                                                                 : std_logic_vector(1 downto 0);   -- rotary_in_s1_translator:av_address -> rotary_in:address
	signal rotary_in_s1_translator_avalon_anti_slave_0_readdata                                                                : std_logic_vector(31 downto 0);  -- rotary_in:readdata -> rotary_in_s1_translator:av_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                                             : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	signal cpu_instruction_master_translator_avalon_universal_master_0_burstcount                                              : std_logic_vector(2 downto 0);   -- cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_instruction_master_translator_avalon_universal_master_0_writedata                                               : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_instruction_master_translator_avalon_universal_master_0_address                                                 : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_instruction_master_translator_avalon_universal_master_0_lock                                                    : std_logic;                      -- cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_instruction_master_translator_avalon_universal_master_0_write                                                   : std_logic;                      -- cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_instruction_master_translator_avalon_universal_master_0_read                                                    : std_logic;                      -- cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdata                                                : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                                             : std_logic;                      -- cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_instruction_master_translator_avalon_universal_master_0_byteenable                                              : std_logic_vector(3 downto 0);   -- cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                                           : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest                           : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_waitrequest
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount                            : std_logic_vector(1 downto 0);   -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_burstcount -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata                             : std_logic_vector(15 downto 0);  -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_writedata -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_address                               : std_logic_vector(31 downto 0);  -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_address -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock                                  : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_lock -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_write                                 : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_write -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_read                                  : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_read -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata                              : std_logic_vector(15 downto 0);  -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_readdata
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess                           : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_debugaccess -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable                            : std_logic_vector(1 downto 0);   -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_byteenable -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid                         : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_readdatavalid
	signal cpu_data_master_translator_avalon_universal_master_0_waitrequest                                                    : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	signal cpu_data_master_translator_avalon_universal_master_0_burstcount                                                     : std_logic_vector(2 downto 0);   -- cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_data_master_translator_avalon_universal_master_0_writedata                                                      : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_data_master_translator_avalon_universal_master_0_address                                                        : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_data_master_translator_avalon_universal_master_0_lock                                                           : std_logic;                      -- cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_data_master_translator_avalon_universal_master_0_write                                                          : std_logic;                      -- cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_data_master_translator_avalon_universal_master_0_read                                                           : std_logic;                      -- cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_data_master_translator_avalon_universal_master_0_readdata                                                       : std_logic_vector(31 downto 0);  -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_debugaccess                                                    : std_logic;                      -- cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_data_master_translator_avalon_universal_master_0_byteenable                                                     : std_logic_vector(3 downto 0);   -- cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_data_master_translator_avalon_universal_master_0_readdatavalid                                                  : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                                      : std_logic;                      -- cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                                       : std_logic_vector(2 downto 0);   -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                                        : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                                          : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                                            : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                                             : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                                             : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                                         : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                    : std_logic;                      -- cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                                      : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                                       : std_logic_vector(3 downto 0);   -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                               : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                                     : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                             : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                                      : std_logic_vector(109 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                                     : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                            : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                  : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                          : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                   : std_logic_vector(109 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                  : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                 : std_logic_vector(33 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                 : std_logic_vector(33 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- SRAM_avalon_sram_slave_translator:uav_waitrequest -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(1 downto 0);   -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SRAM_avalon_sram_slave_translator:uav_burstcount
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(15 downto 0);  -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SRAM_avalon_sram_slave_translator:uav_writedata
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(31 downto 0);  -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> SRAM_avalon_sram_slave_translator:uav_address
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> SRAM_avalon_sram_slave_translator:uav_write
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SRAM_avalon_sram_slave_translator:uav_lock
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> SRAM_avalon_sram_slave_translator:uav_read
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(15 downto 0);  -- SRAM_avalon_sram_slave_translator:uav_readdata -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- SRAM_avalon_sram_slave_translator:uav_readdatavalid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SRAM_avalon_sram_slave_translator:uav_debugaccess
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(1 downto 0);   -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SRAM_avalon_sram_slave_translator:uav_byteenable
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(91 downto 0);  -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(91 downto 0);  -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(17 downto 0);  -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                               : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                : std_logic_vector(17 downto 0);  -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                               : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(109 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(109 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                           : std_logic_vector(33 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                           : std_logic;                      -- sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                            : std_logic_vector(2 downto 0);   -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                             : std_logic_vector(31 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address                                               : std_logic_vector(31 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write                                                 : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                  : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read                                                  : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                              : std_logic_vector(31 downto 0);  -- sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                         : std_logic;                      -- sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                           : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                            : std_logic_vector(3 downto 0);   -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                    : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                          : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                  : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                           : std_logic_vector(109 downto 0); -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                          : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                 : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                       : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                               : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                        : std_logic_vector(109 downto 0); -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                       : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                      : std_logic_vector(33 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                      : std_logic_vector(33 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                        : std_logic;                      -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                         : std_logic_vector(2 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                          : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                            : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                           : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                      : std_logic;                      -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                         : std_logic_vector(3 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                 : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                       : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                        : std_logic_vector(109 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                       : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                            : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                     : std_logic_vector(109 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                   : std_logic_vector(33 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                   : std_logic_vector(33 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                             : std_logic;                      -- red_led_pio_s1_translator:uav_waitrequest -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                              : std_logic_vector(2 downto 0);   -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> red_led_pio_s1_translator:uav_burstcount
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                               : std_logic_vector(31 downto 0);  -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> red_led_pio_s1_translator:uav_writedata
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address                                                 : std_logic_vector(31 downto 0);  -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> red_led_pio_s1_translator:uav_address
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write                                                   : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> red_led_pio_s1_translator:uav_write
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                    : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> red_led_pio_s1_translator:uav_lock
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read                                                    : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> red_led_pio_s1_translator:uav_read
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                : std_logic_vector(31 downto 0);  -- red_led_pio_s1_translator:uav_readdata -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                           : std_logic;                      -- red_led_pio_s1_translator:uav_readdatavalid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                             : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> red_led_pio_s1_translator:uav_debugaccess
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                              : std_logic_vector(3 downto 0);   -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> red_led_pio_s1_translator:uav_byteenable
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                      : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                            : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                    : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                             : std_logic_vector(109 downto 0); -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                            : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                   : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                         : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                 : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                          : std_logic_vector(109 downto 0); -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                         : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                       : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                        : std_logic_vector(33 downto 0);  -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                       : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                       : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                        : std_logic_vector(33 downto 0);  -- red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                       : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator:uav_waitrequest -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_burstcount
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_writedata
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(31 downto 0);  -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_address
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_write
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_lock
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_read
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- VGA_Character_buffer_avalon_char_control_slave_translator:uav_readdata -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator:uav_readdatavalid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_debugaccess
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_byteenable
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(109 downto 0); -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(109 downto 0); -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid       : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data        : std_logic_vector(33 downto 0);  -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready       : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_waitrequest -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(0 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_burstcount
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(7 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_writedata
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(31 downto 0);  -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_address
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_write
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_lock
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_read
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(7 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_readdata -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_readdatavalid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_debugaccess
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(0 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_byteenable
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(82 downto 0);  -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(82 downto 0);  -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(9 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid        : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data         : std_logic_vector(9 downto 0);   -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready        : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator:uav_waitrequest -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);   -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_burstcount
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0);  -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_writedata
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(31 downto 0);  -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_address
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_write
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_lock
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_read
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0);  -- VGA_Pixel_Buffer_avalon_control_slave_translator:uav_readdata -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator:uav_readdatavalid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_debugaccess
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);   -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_byteenable
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(109 downto 0); -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(109 downto 0); -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(33 downto 0);  -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                 : std_logic_vector(33 downto 0);  -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                           : std_logic;                      -- green_led_pio_s1_translator:uav_waitrequest -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                            : std_logic_vector(2 downto 0);   -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> green_led_pio_s1_translator:uav_burstcount
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                             : std_logic_vector(31 downto 0);  -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> green_led_pio_s1_translator:uav_writedata
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address                                               : std_logic_vector(31 downto 0);  -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> green_led_pio_s1_translator:uav_address
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write                                                 : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> green_led_pio_s1_translator:uav_write
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                  : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> green_led_pio_s1_translator:uav_lock
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read                                                  : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> green_led_pio_s1_translator:uav_read
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                              : std_logic_vector(31 downto 0);  -- green_led_pio_s1_translator:uav_readdata -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                         : std_logic;                      -- green_led_pio_s1_translator:uav_readdatavalid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                           : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> green_led_pio_s1_translator:uav_debugaccess
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                            : std_logic_vector(3 downto 0);   -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> green_led_pio_s1_translator:uav_byteenable
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                    : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                          : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                  : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                           : std_logic_vector(109 downto 0); -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                          : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                 : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                       : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                               : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                        : std_logic_vector(109 downto 0); -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                       : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                     : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                      : std_logic_vector(33 downto 0);  -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                     : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                     : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                      : std_logic_vector(33 downto 0);  -- green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                     : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                              : std_logic;                      -- control_in_s1_translator:uav_waitrequest -> control_in_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                               : std_logic_vector(2 downto 0);   -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> control_in_s1_translator:uav_burstcount
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                : std_logic_vector(31 downto 0);  -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> control_in_s1_translator:uav_writedata
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_address                                                  : std_logic_vector(31 downto 0);  -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_address -> control_in_s1_translator:uav_address
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_write                                                    : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_write -> control_in_s1_translator:uav_write
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                     : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_lock -> control_in_s1_translator:uav_lock
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_read                                                     : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_read -> control_in_s1_translator:uav_read
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                 : std_logic_vector(31 downto 0);  -- control_in_s1_translator:uav_readdata -> control_in_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                            : std_logic;                      -- control_in_s1_translator:uav_readdatavalid -> control_in_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                              : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> control_in_s1_translator:uav_debugaccess
	signal control_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                               : std_logic_vector(3 downto 0);   -- control_in_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> control_in_s1_translator:uav_byteenable
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                       : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                             : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                     : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                              : std_logic_vector(109 downto 0); -- control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                             : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                    : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                          : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                  : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                           : std_logic_vector(109 downto 0); -- control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                          : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                        : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                         : std_logic_vector(33 downto 0);  -- control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                        : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                        : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                         : std_logic_vector(33 downto 0);  -- control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                        : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                             : std_logic;                      -- control_out_s1_translator:uav_waitrequest -> control_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                              : std_logic_vector(2 downto 0);   -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> control_out_s1_translator:uav_burstcount
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                               : std_logic_vector(31 downto 0);  -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> control_out_s1_translator:uav_writedata
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_address                                                 : std_logic_vector(31 downto 0);  -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> control_out_s1_translator:uav_address
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_write                                                   : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> control_out_s1_translator:uav_write
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                    : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> control_out_s1_translator:uav_lock
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_read                                                    : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> control_out_s1_translator:uav_read
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                : std_logic_vector(31 downto 0);  -- control_out_s1_translator:uav_readdata -> control_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                           : std_logic;                      -- control_out_s1_translator:uav_readdatavalid -> control_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                             : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> control_out_s1_translator:uav_debugaccess
	signal control_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                              : std_logic_vector(3 downto 0);   -- control_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> control_out_s1_translator:uav_byteenable
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                      : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                            : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                    : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                             : std_logic_vector(109 downto 0); -- control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                            : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                   : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                         : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                 : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                          : std_logic_vector(109 downto 0); -- control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                         : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                       : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                        : std_logic_vector(33 downto 0);  -- control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                       : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                       : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                        : std_logic_vector(33 downto 0);  -- control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                       : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                : std_logic;                      -- FFT_in_0_s1_translator:uav_waitrequest -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                 : std_logic_vector(2 downto 0);   -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_0_s1_translator:uav_burstcount
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                  : std_logic_vector(31 downto 0);  -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_0_s1_translator:uav_writedata
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                                    : std_logic_vector(31 downto 0);  -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_0_s1_translator:uav_address
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                                      : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_0_s1_translator:uav_write
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                       : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_0_s1_translator:uav_lock
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                                       : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_0_s1_translator:uav_read
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                   : std_logic_vector(31 downto 0);  -- FFT_in_0_s1_translator:uav_readdata -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                              : std_logic;                      -- FFT_in_0_s1_translator:uav_readdatavalid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_0_s1_translator:uav_debugaccess
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                 : std_logic_vector(3 downto 0);   -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_0_s1_translator:uav_byteenable
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                         : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                               : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                       : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                : std_logic_vector(109 downto 0); -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                               : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                      : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                            : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                    : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                             : std_logic_vector(109 downto 0); -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                            : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                          : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                          : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                          : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                          : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                : std_logic;                      -- FFT_in_1_s1_translator:uav_waitrequest -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                 : std_logic_vector(2 downto 0);   -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_1_s1_translator:uav_burstcount
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                  : std_logic_vector(31 downto 0);  -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_1_s1_translator:uav_writedata
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_address                                                    : std_logic_vector(31 downto 0);  -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_1_s1_translator:uav_address
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_write                                                      : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_1_s1_translator:uav_write
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                       : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_1_s1_translator:uav_lock
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_read                                                       : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_1_s1_translator:uav_read
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                   : std_logic_vector(31 downto 0);  -- FFT_in_1_s1_translator:uav_readdata -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                              : std_logic;                      -- FFT_in_1_s1_translator:uav_readdatavalid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_1_s1_translator:uav_debugaccess
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                 : std_logic_vector(3 downto 0);   -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_1_s1_translator:uav_byteenable
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                         : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                               : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                       : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                : std_logic_vector(109 downto 0); -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                               : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                      : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                            : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                    : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                             : std_logic_vector(109 downto 0); -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                            : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                          : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                          : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                          : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                          : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                : std_logic;                      -- FFT_in_2_s1_translator:uav_waitrequest -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                 : std_logic_vector(2 downto 0);   -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_2_s1_translator:uav_burstcount
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                  : std_logic_vector(31 downto 0);  -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_2_s1_translator:uav_writedata
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_address                                                    : std_logic_vector(31 downto 0);  -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_2_s1_translator:uav_address
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_write                                                      : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_2_s1_translator:uav_write
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                       : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_2_s1_translator:uav_lock
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_read                                                       : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_2_s1_translator:uav_read
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                   : std_logic_vector(31 downto 0);  -- FFT_in_2_s1_translator:uav_readdata -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                              : std_logic;                      -- FFT_in_2_s1_translator:uav_readdatavalid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_2_s1_translator:uav_debugaccess
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                 : std_logic_vector(3 downto 0);   -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_2_s1_translator:uav_byteenable
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                         : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                               : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                       : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                : std_logic_vector(109 downto 0); -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                               : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                      : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                            : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                    : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                             : std_logic_vector(109 downto 0); -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                            : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                          : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                          : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                          : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                          : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                : std_logic;                      -- FFT_in_3_s1_translator:uav_waitrequest -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                 : std_logic_vector(2 downto 0);   -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_3_s1_translator:uav_burstcount
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                  : std_logic_vector(31 downto 0);  -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_3_s1_translator:uav_writedata
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_address                                                    : std_logic_vector(31 downto 0);  -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_3_s1_translator:uav_address
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_write                                                      : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_3_s1_translator:uav_write
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                       : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_3_s1_translator:uav_lock
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_read                                                       : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_3_s1_translator:uav_read
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                   : std_logic_vector(31 downto 0);  -- FFT_in_3_s1_translator:uav_readdata -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                              : std_logic;                      -- FFT_in_3_s1_translator:uav_readdatavalid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_3_s1_translator:uav_debugaccess
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                 : std_logic_vector(3 downto 0);   -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_3_s1_translator:uav_byteenable
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                         : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                               : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                       : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                : std_logic_vector(109 downto 0); -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                               : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                      : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                            : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                    : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                             : std_logic_vector(109 downto 0); -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                            : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                          : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                          : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                          : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                           : std_logic_vector(33 downto 0);  -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                          : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                               : std_logic;                      -- rotary_in_s1_translator:uav_waitrequest -> rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                : std_logic_vector(2 downto 0);   -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> rotary_in_s1_translator:uav_burstcount
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                 : std_logic_vector(31 downto 0);  -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> rotary_in_s1_translator:uav_writedata
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_address                                                   : std_logic_vector(31 downto 0);  -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_address -> rotary_in_s1_translator:uav_address
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_write                                                     : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_write -> rotary_in_s1_translator:uav_write
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                      : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_lock -> rotary_in_s1_translator:uav_lock
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_read                                                      : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_read -> rotary_in_s1_translator:uav_read
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                  : std_logic_vector(31 downto 0);  -- rotary_in_s1_translator:uav_readdata -> rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                             : std_logic;                      -- rotary_in_s1_translator:uav_readdatavalid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                               : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rotary_in_s1_translator:uav_debugaccess
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                : std_logic_vector(3 downto 0);   -- rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> rotary_in_s1_translator:uav_byteenable
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                        : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                              : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                      : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                               : std_logic_vector(109 downto 0); -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                              : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                     : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                           : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                   : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                            : std_logic_vector(109 downto 0); -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                           : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                         : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                          : std_logic_vector(33 downto 0);  -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                         : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                         : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                          : std_logic_vector(33 downto 0);  -- rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                         : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                                    : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                                          : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                                  : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                                           : std_logic_vector(108 downto 0); -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                                          : std_logic;                      -- addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket                  : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid                        : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket                : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data                         : std_logic_vector(90 downto 0);  -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready                        : std_logic;                      -- addr_router_001:sink_ready -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                                           : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                                                 : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                                         : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                                                  : std_logic_vector(108 downto 0); -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                                                 : std_logic;                      -- addr_router_002:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                                      : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                                            : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                                    : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                                             : std_logic_vector(108 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                                            : std_logic;                      -- id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(90 downto 0);  -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_001:sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(108 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                      -- id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                           : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                 : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                         : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data                                                  : std_logic_vector(108 downto 0); -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                 : std_logic;                      -- id_router_003:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                               : std_logic_vector(108 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                              : std_logic;                      -- id_router_004:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                             : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                   : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                           : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data                                                    : std_logic_vector(108 downto 0); -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                   : std_logic;                      -- id_router_005:sink_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(108 downto 0); -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_006:sink_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(81 downto 0);  -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                      -- id_router_007:sink_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(108 downto 0); -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                      -- id_router_008:sink_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                           : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                 : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                         : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data                                                  : std_logic_vector(108 downto 0); -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                 : std_logic;                      -- id_router_009:sink_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                              : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                    : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                            : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rp_data                                                     : std_logic_vector(108 downto 0); -- control_in_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal control_in_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                    : std_logic;                      -- id_router_010:sink_ready -> control_in_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                             : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                   : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                           : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rp_data                                                    : std_logic_vector(108 downto 0); -- control_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal control_out_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                   : std_logic;                      -- id_router_011:sink_ready -> control_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                      : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                              : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                                       : std_logic_vector(108 downto 0); -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                      : std_logic;                      -- id_router_012:sink_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                      : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                              : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_data                                                       : std_logic_vector(108 downto 0); -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                      : std_logic;                      -- id_router_013:sink_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                      : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                              : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_data                                                       : std_logic_vector(108 downto 0); -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                      : std_logic;                      -- id_router_014:sink_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                      : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                              : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_data                                                       : std_logic_vector(108 downto 0); -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	signal fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                      : std_logic;                      -- id_router_015:sink_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                               : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                     : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                             : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_data                                                      : std_logic_vector(108 downto 0); -- rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	signal rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                     : std_logic;                      -- id_router_016:sink_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal burst_adapter_source0_endofpacket                                                                                   : std_logic;                      -- burst_adapter:source0_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                                         : std_logic;                      -- burst_adapter:source0_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                                 : std_logic;                      -- burst_adapter:source0_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                                          : std_logic_vector(90 downto 0);  -- burst_adapter:source0_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                                         : std_logic;                      -- SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                                       : std_logic_vector(16 downto 0);  -- burst_adapter:source0_channel -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                                               : std_logic;                      -- burst_adapter_001:source0_endofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                                     : std_logic;                      -- burst_adapter_001:source0_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                                             : std_logic;                      -- burst_adapter_001:source0_startofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                                      : std_logic_vector(81 downto 0);  -- burst_adapter_001:source0_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                                     : std_logic;                      -- VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                                   : std_logic_vector(16 downto 0);  -- burst_adapter_001:source0_channel -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                                      : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux:reset, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:in_reset, crosser_007:out_reset, crosser_008:out_reset, crosser_009:out_reset, id_router:reset, id_router_002:reset, irq_mapper:reset, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_002:reset, rsp_xbar_mux:reset, rsp_xbar_mux_002:reset, rst_controller_reset_out_reset:in, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset]
	signal external_clocks_sys_clk_reset_reset                                                                                 : std_logic;                      -- external_clocks:sys_reset_n -> external_clocks_sys_clk_reset_reset:in
	signal rst_controller_001_reset_out_reset                                                                                  : std_logic;                      -- rst_controller_001:reset_out -> [FFT_in_0_s1_translator:reset, FFT_in_0_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_1_s1_translator:reset, FFT_in_1_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_2_s1_translator:reset, FFT_in_2_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_3_s1_translator:reset, FFT_in_3_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, control_in_s1_translator:reset, control_in_s1_translator_avalon_universal_slave_0_agent:reset, control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, control_out_s1_translator:reset, control_out_s1_translator_avalon_universal_slave_0_agent:reset, control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, external_clocks:reset, green_led_pio_s1_translator:reset, green_led_pio_s1_translator_avalon_universal_slave_0_agent:reset, green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, red_led_pio_s1_translator:reset, red_led_pio_s1_translator_avalon_universal_slave_0_agent:reset, red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rotary_in_s1_translator:reset, rotary_in_s1_translator_avalon_universal_slave_0_agent:reset, rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rst_controller_001_reset_out_reset:in, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal rst_controller_002_reset_out_reset                                                                                  : std_logic;                      -- rst_controller_002:reset_out -> [Alpha_Blending:reset, SRAM:reset, SRAM_avalon_sram_slave_translator:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Character_buffer:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Character_buffer_avalon_char_control_slave_translator:reset, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Dual_Clock_FIFO:reset_stream_in, VGA_Pixel_Buffer:reset, VGA_Pixel_Buffer_avalon_control_slave_translator:reset, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:reset, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, VGA_Scaler:reset, VGA_pixel_RGB_Resampler:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux_001:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:in_reset, crosser_008:in_reset, crosser_009:in_reset, id_router_001:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset]
	signal cpu_jtag_debug_module_reset_reset                                                                                   : std_logic;                      -- cpu:jtag_debug_module_resetrequest -> [rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	signal rst_controller_003_reset_out_reset                                                                                  : std_logic;                      -- rst_controller_003:reset_out -> [VGA_Controller:reset, VGA_Dual_Clock_FIFO:reset_stream_out]
	signal cmd_xbar_demux_src0_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                                           : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                                            : std_logic_vector(108 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                                         : std_logic_vector(16 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                                           : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                                        : std_logic_vector(90 downto 0);  -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                                       : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_002_src0_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_002_src0_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_002_src0_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_002_src0_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_002_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_002_src0_ready                                                                                       : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_002:src0_ready
	signal cmd_xbar_demux_002_src2_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src2_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src2_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src2_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src2_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src3_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src3_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src3_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src3_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src3_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src3_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src3_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src3_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src3_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src3_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src4_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src4_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src4_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src4_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src4_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src4_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src4_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src4_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src4_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src4_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src5_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src5_endofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src5_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src5_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src5_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src5_startofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src5_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src5_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src5_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src5_channel -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src9_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src9_endofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src9_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src9_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src9_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src9_startofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src9_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src9_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src9_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src9_channel -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src10_endofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_002:src10_endofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src10_valid                                                                                      : std_logic;                      -- cmd_xbar_demux_002:src10_valid -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src10_startofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_002:src10_startofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src10_data                                                                                       : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src10_data -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src10_channel                                                                                    : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src10_channel -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src11_endofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_002:src11_endofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src11_valid                                                                                      : std_logic;                      -- cmd_xbar_demux_002:src11_valid -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src11_startofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_002:src11_startofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src11_data                                                                                       : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src11_data -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src11_channel                                                                                    : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src11_channel -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src12_endofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_002:src12_endofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src12_valid                                                                                      : std_logic;                      -- cmd_xbar_demux_002:src12_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src12_startofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_002:src12_startofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src12_data                                                                                       : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src12_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src12_channel                                                                                    : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src12_channel -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src13_endofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_002:src13_endofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src13_valid                                                                                      : std_logic;                      -- cmd_xbar_demux_002:src13_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src13_startofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_002:src13_startofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src13_data                                                                                       : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src13_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src13_channel                                                                                    : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src13_channel -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src14_endofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_002:src14_endofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src14_valid                                                                                      : std_logic;                      -- cmd_xbar_demux_002:src14_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src14_startofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_002:src14_startofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src14_data                                                                                       : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src14_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src14_channel                                                                                    : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src14_channel -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src15_endofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_002:src15_endofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src15_valid                                                                                      : std_logic;                      -- cmd_xbar_demux_002:src15_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src15_startofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_002:src15_startofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src15_data                                                                                       : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src15_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src15_channel                                                                                    : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src15_channel -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src16_endofpacket                                                                                : std_logic;                      -- cmd_xbar_demux_002:src16_endofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_002_src16_valid                                                                                      : std_logic;                      -- cmd_xbar_demux_002:src16_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_002_src16_startofpacket                                                                              : std_logic;                      -- cmd_xbar_demux_002:src16_startofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_002_src16_data                                                                                       : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src16_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_002_src16_channel                                                                                    : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src16_channel -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                                     : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                                           : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                                   : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                                            : std_logic_vector(108 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                                         : std_logic_vector(16 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                                           : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                                     : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                                           : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_002:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                                   : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                                            : std_logic_vector(108 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_002:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                                         : std_logic_vector(16 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_002:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                                           : std_logic;                      -- rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                                        : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_001:src1_data -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_001_src1_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_001:src1_channel -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_002_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_002:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_002:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_002:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_002:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_002:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_002:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_002:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_002:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_002:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_002:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_002:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_002:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_002:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_002:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_002:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_002:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_002:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_002:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_002:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_002:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_002:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_002:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_002:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_002:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_002:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_002:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_002:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_002:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_002:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_002:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_002:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_002:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_002:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_002:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_002:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_002:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_002:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_002:sink14_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_002:sink14_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_002:sink14_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_002:sink14_data
	signal rsp_xbar_demux_014_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_002:sink14_channel
	signal rsp_xbar_demux_014_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink14_ready -> rsp_xbar_demux_014:src0_ready
	signal rsp_xbar_demux_015_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_002:sink15_endofpacket
	signal rsp_xbar_demux_015_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_002:sink15_valid
	signal rsp_xbar_demux_015_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_002:sink15_startofpacket
	signal rsp_xbar_demux_015_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_002:sink15_data
	signal rsp_xbar_demux_015_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_002:sink15_channel
	signal rsp_xbar_demux_015_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink15_ready -> rsp_xbar_demux_015:src0_ready
	signal rsp_xbar_demux_016_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_002:sink16_endofpacket
	signal rsp_xbar_demux_016_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_002:sink16_valid
	signal rsp_xbar_demux_016_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_002:sink16_startofpacket
	signal rsp_xbar_demux_016_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_002:sink16_data
	signal rsp_xbar_demux_016_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_002:sink16_channel
	signal rsp_xbar_demux_016_src0_ready                                                                                       : std_logic;                      -- rsp_xbar_mux_002:sink16_ready -> rsp_xbar_demux_016:src0_ready
	signal addr_router_src_endofpacket                                                                                         : std_logic;                      -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                                               : std_logic;                      -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                                       : std_logic;                      -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                                : std_logic_vector(108 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                                             : std_logic_vector(16 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                                               : std_logic;                      -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                                        : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                              : std_logic;                      -- rsp_xbar_mux:src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                                      : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                                               : std_logic_vector(108 downto 0); -- rsp_xbar_mux:src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                                            : std_logic_vector(16 downto 0);  -- rsp_xbar_mux:src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                                              : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                                     : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                                           : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                                   : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                                            : std_logic_vector(90 downto 0);  -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                                         : std_logic_vector(16 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                                           : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_demux_001_src1_ready                                                                                       : std_logic;                      -- VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src1_ready
	signal addr_router_002_src_endofpacket                                                                                     : std_logic;                      -- addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	signal addr_router_002_src_valid                                                                                           : std_logic;                      -- addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	signal addr_router_002_src_startofpacket                                                                                   : std_logic;                      -- addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	signal addr_router_002_src_data                                                                                            : std_logic_vector(108 downto 0); -- addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	signal addr_router_002_src_channel                                                                                         : std_logic_vector(16 downto 0);  -- addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	signal addr_router_002_src_ready                                                                                           : std_logic;                      -- cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	signal rsp_xbar_mux_002_src_endofpacket                                                                                    : std_logic;                      -- rsp_xbar_mux_002:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_002_src_valid                                                                                          : std_logic;                      -- rsp_xbar_mux_002:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_002_src_startofpacket                                                                                  : std_logic;                      -- rsp_xbar_mux_002:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_002_src_data                                                                                           : std_logic_vector(108 downto 0); -- rsp_xbar_mux_002:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_002_src_channel                                                                                        : std_logic_vector(16 downto 0);  -- rsp_xbar_mux_002:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_002_src_ready                                                                                          : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                                        : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                              : std_logic;                      -- cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                                      : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                               : std_logic_vector(108 downto 0); -- cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                                            : std_logic_vector(16 downto 0);  -- cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                              : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                                           : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                                 : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                                         : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                                  : std_logic_vector(108 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                               : std_logic_vector(16 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                                 : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                                    : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> burst_adapter:sink0_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                                          : std_logic;                      -- cmd_xbar_mux_001:src_valid -> burst_adapter:sink0_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                                  : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> burst_adapter:sink0_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                                           : std_logic_vector(90 downto 0);  -- cmd_xbar_mux_001:src_data -> burst_adapter:sink0_data
	signal cmd_xbar_mux_001_src_channel                                                                                        : std_logic_vector(16 downto 0);  -- cmd_xbar_mux_001:src_channel -> burst_adapter:sink0_channel
	signal cmd_xbar_mux_001_src_ready                                                                                          : std_logic;                      -- burst_adapter:sink0_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                                       : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                                             : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                                     : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                                              : std_logic_vector(90 downto 0);  -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_demux_002_src2_ready                                                                                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src2_ready
	signal id_router_002_src_endofpacket                                                                                       : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                                             : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                                     : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_demux_002_src3_ready                                                                                       : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src3_ready
	signal id_router_003_src_endofpacket                                                                                       : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                                             : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                                     : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_002_src4_ready                                                                                       : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src4_ready
	signal id_router_004_src_endofpacket                                                                                       : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                             : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                                     : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_002_src5_ready                                                                                       : std_logic;                      -- red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src5_ready
	signal id_router_005_src_endofpacket                                                                                       : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                             : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                                     : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal crosser_out_ready                                                                                                   : std_logic;                      -- VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	signal id_router_006_src_endofpacket                                                                                       : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                             : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                                     : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal crosser_006_out_ready                                                                                               : std_logic;                      -- burst_adapter_001:sink0_ready -> crosser_006:out_ready
	signal id_router_007_src_endofpacket                                                                                       : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                             : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                                     : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                              : std_logic_vector(81 downto 0);  -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal crosser_001_out_ready                                                                                               : std_logic;                      -- VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	signal id_router_008_src_endofpacket                                                                                       : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                                             : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                                     : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_002_src9_ready                                                                                       : std_logic;                      -- green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src9_ready
	signal id_router_009_src_endofpacket                                                                                       : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                                             : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                                     : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_002_src10_ready                                                                                      : std_logic;                      -- control_in_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src10_ready
	signal id_router_010_src_endofpacket                                                                                       : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                                             : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                                     : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_002_src11_ready                                                                                      : std_logic;                      -- control_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src11_ready
	signal id_router_011_src_endofpacket                                                                                       : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                                             : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                                     : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_002_src12_ready                                                                                      : std_logic;                      -- FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src12_ready
	signal id_router_012_src_endofpacket                                                                                       : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                                             : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                                     : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_demux_002_src13_ready                                                                                      : std_logic;                      -- FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src13_ready
	signal id_router_013_src_endofpacket                                                                                       : std_logic;                      -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                                             : std_logic;                      -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                                                     : std_logic;                      -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal cmd_xbar_demux_002_src14_ready                                                                                      : std_logic;                      -- FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src14_ready
	signal id_router_014_src_endofpacket                                                                                       : std_logic;                      -- id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal id_router_014_src_valid                                                                                             : std_logic;                      -- id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	signal id_router_014_src_startofpacket                                                                                     : std_logic;                      -- id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal id_router_014_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	signal id_router_014_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	signal id_router_014_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	signal cmd_xbar_demux_002_src15_ready                                                                                      : std_logic;                      -- FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src15_ready
	signal id_router_015_src_endofpacket                                                                                       : std_logic;                      -- id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	signal id_router_015_src_valid                                                                                             : std_logic;                      -- id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	signal id_router_015_src_startofpacket                                                                                     : std_logic;                      -- id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	signal id_router_015_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	signal id_router_015_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	signal id_router_015_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	signal cmd_xbar_demux_002_src16_ready                                                                                      : std_logic;                      -- rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src16_ready
	signal id_router_016_src_endofpacket                                                                                       : std_logic;                      -- id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	signal id_router_016_src_valid                                                                                             : std_logic;                      -- id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	signal id_router_016_src_startofpacket                                                                                     : std_logic;                      -- id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	signal id_router_016_src_data                                                                                              : std_logic_vector(108 downto 0); -- id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	signal id_router_016_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	signal id_router_016_src_ready                                                                                             : std_logic;                      -- rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                                     : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                                           : std_logic;                      -- cmd_xbar_demux:src1_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                                   : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_src1_data                                                                                            : std_logic_vector(108 downto 0); -- cmd_xbar_demux:src1_data -> width_adapter:in_data
	signal cmd_xbar_demux_src1_channel                                                                                         : std_logic_vector(16 downto 0);  -- cmd_xbar_demux:src1_channel -> width_adapter:in_channel
	signal cmd_xbar_demux_src1_ready                                                                                           : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_002_src1_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src1_endofpacket -> width_adapter_001:in_endofpacket
	signal cmd_xbar_demux_002_src1_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src1_valid -> width_adapter_001:in_valid
	signal cmd_xbar_demux_002_src1_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src1_startofpacket -> width_adapter_001:in_startofpacket
	signal cmd_xbar_demux_002_src1_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src1_data -> width_adapter_001:in_data
	signal cmd_xbar_demux_002_src1_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src1_channel -> width_adapter_001:in_channel
	signal cmd_xbar_demux_002_src1_ready                                                                                       : std_logic;                      -- width_adapter_001:in_ready -> cmd_xbar_demux_002:src1_ready
	signal cmd_xbar_demux_002_src7_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src7_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_demux_002_src7_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src7_valid -> width_adapter_002:in_valid
	signal cmd_xbar_demux_002_src7_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src7_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_demux_002_src7_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src7_data -> width_adapter_002:in_data
	signal cmd_xbar_demux_002_src7_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src7_channel -> width_adapter_002:in_channel
	signal cmd_xbar_demux_002_src7_ready                                                                                       : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_demux_002:src7_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> width_adapter_003:in_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> width_adapter_003:in_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> width_adapter_003:in_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                                        : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_001:src0_data -> width_adapter_003:in_data
	signal rsp_xbar_demux_001_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_001:src0_channel -> width_adapter_003:in_channel
	signal rsp_xbar_demux_001_src0_ready                                                                                       : std_logic;                      -- width_adapter_003:in_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src2_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_001:src2_endofpacket -> width_adapter_004:in_endofpacket
	signal rsp_xbar_demux_001_src2_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_001:src2_valid -> width_adapter_004:in_valid
	signal rsp_xbar_demux_001_src2_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_001:src2_startofpacket -> width_adapter_004:in_startofpacket
	signal rsp_xbar_demux_001_src2_data                                                                                        : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_001:src2_data -> width_adapter_004:in_data
	signal rsp_xbar_demux_001_src2_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_001:src2_channel -> width_adapter_004:in_channel
	signal rsp_xbar_demux_001_src2_ready                                                                                       : std_logic;                      -- width_adapter_004:in_ready -> rsp_xbar_demux_001:src2_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> width_adapter_005:in_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> width_adapter_005:in_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> width_adapter_005:in_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                                        : std_logic_vector(81 downto 0);  -- rsp_xbar_demux_007:src0_data -> width_adapter_005:in_data
	signal rsp_xbar_demux_007_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_007:src0_channel -> width_adapter_005:in_channel
	signal rsp_xbar_demux_007_src0_ready                                                                                       : std_logic;                      -- width_adapter_005:in_ready -> rsp_xbar_demux_007:src0_ready
	signal crosser_out_endofpacket                                                                                             : std_logic;                      -- crosser:out_endofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal crosser_out_valid                                                                                                   : std_logic;                      -- crosser:out_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal crosser_out_startofpacket                                                                                           : std_logic;                      -- crosser:out_startofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal crosser_out_data                                                                                                    : std_logic_vector(108 downto 0); -- crosser:out_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal crosser_out_channel                                                                                                 : std_logic_vector(16 downto 0);  -- crosser:out_channel -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src6_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src6_endofpacket -> crosser:in_endofpacket
	signal cmd_xbar_demux_002_src6_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src6_valid -> crosser:in_valid
	signal cmd_xbar_demux_002_src6_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src6_startofpacket -> crosser:in_startofpacket
	signal cmd_xbar_demux_002_src6_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src6_data -> crosser:in_data
	signal cmd_xbar_demux_002_src6_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src6_channel -> crosser:in_channel
	signal cmd_xbar_demux_002_src6_ready                                                                                       : std_logic;                      -- crosser:in_ready -> cmd_xbar_demux_002:src6_ready
	signal crosser_001_out_endofpacket                                                                                         : std_logic;                      -- crosser_001:out_endofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal crosser_001_out_valid                                                                                               : std_logic;                      -- crosser_001:out_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal crosser_001_out_startofpacket                                                                                       : std_logic;                      -- crosser_001:out_startofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal crosser_001_out_data                                                                                                : std_logic_vector(108 downto 0); -- crosser_001:out_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal crosser_001_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_001:out_channel -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_002_src8_endofpacket                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src8_endofpacket -> crosser_001:in_endofpacket
	signal cmd_xbar_demux_002_src8_valid                                                                                       : std_logic;                      -- cmd_xbar_demux_002:src8_valid -> crosser_001:in_valid
	signal cmd_xbar_demux_002_src8_startofpacket                                                                               : std_logic;                      -- cmd_xbar_demux_002:src8_startofpacket -> crosser_001:in_startofpacket
	signal cmd_xbar_demux_002_src8_data                                                                                        : std_logic_vector(108 downto 0); -- cmd_xbar_demux_002:src8_data -> crosser_001:in_data
	signal cmd_xbar_demux_002_src8_channel                                                                                     : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src8_channel -> crosser_001:in_channel
	signal cmd_xbar_demux_002_src8_ready                                                                                       : std_logic;                      -- crosser_001:in_ready -> cmd_xbar_demux_002:src8_ready
	signal crosser_002_out_endofpacket                                                                                         : std_logic;                      -- crosser_002:out_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	signal crosser_002_out_valid                                                                                               : std_logic;                      -- crosser_002:out_valid -> rsp_xbar_mux_002:sink6_valid
	signal crosser_002_out_startofpacket                                                                                       : std_logic;                      -- crosser_002:out_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	signal crosser_002_out_data                                                                                                : std_logic_vector(108 downto 0); -- crosser_002:out_data -> rsp_xbar_mux_002:sink6_data
	signal crosser_002_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_002:out_channel -> rsp_xbar_mux_002:sink6_channel
	signal crosser_002_out_ready                                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink6_ready -> crosser_002:out_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> crosser_002:in_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> crosser_002:in_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> crosser_002:in_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_006:src0_data -> crosser_002:in_data
	signal rsp_xbar_demux_006_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_006:src0_channel -> crosser_002:in_channel
	signal rsp_xbar_demux_006_src0_ready                                                                                       : std_logic;                      -- crosser_002:in_ready -> rsp_xbar_demux_006:src0_ready
	signal crosser_003_out_endofpacket                                                                                         : std_logic;                      -- crosser_003:out_endofpacket -> rsp_xbar_mux_002:sink8_endofpacket
	signal crosser_003_out_valid                                                                                               : std_logic;                      -- crosser_003:out_valid -> rsp_xbar_mux_002:sink8_valid
	signal crosser_003_out_startofpacket                                                                                       : std_logic;                      -- crosser_003:out_startofpacket -> rsp_xbar_mux_002:sink8_startofpacket
	signal crosser_003_out_data                                                                                                : std_logic_vector(108 downto 0); -- crosser_003:out_data -> rsp_xbar_mux_002:sink8_data
	signal crosser_003_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_003:out_channel -> rsp_xbar_mux_002:sink8_channel
	signal crosser_003_out_ready                                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink8_ready -> crosser_003:out_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                                 : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> crosser_003:in_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                                       : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> crosser_003:in_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                               : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> crosser_003:in_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                                        : std_logic_vector(108 downto 0); -- rsp_xbar_demux_008:src0_data -> crosser_003:in_data
	signal rsp_xbar_demux_008_src0_channel                                                                                     : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_008:src0_channel -> crosser_003:in_channel
	signal rsp_xbar_demux_008_src0_ready                                                                                       : std_logic;                      -- crosser_003:in_ready -> rsp_xbar_demux_008:src0_ready
	signal crosser_004_out_endofpacket                                                                                         : std_logic;                      -- crosser_004:out_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal crosser_004_out_valid                                                                                               : std_logic;                      -- crosser_004:out_valid -> cmd_xbar_mux_001:sink0_valid
	signal crosser_004_out_startofpacket                                                                                       : std_logic;                      -- crosser_004:out_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal crosser_004_out_data                                                                                                : std_logic_vector(90 downto 0);  -- crosser_004:out_data -> cmd_xbar_mux_001:sink0_data
	signal crosser_004_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_004:out_channel -> cmd_xbar_mux_001:sink0_channel
	signal crosser_004_out_ready                                                                                               : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> crosser_004:out_ready
	signal width_adapter_src_endofpacket                                                                                       : std_logic;                      -- width_adapter:out_endofpacket -> crosser_004:in_endofpacket
	signal width_adapter_src_valid                                                                                             : std_logic;                      -- width_adapter:out_valid -> crosser_004:in_valid
	signal width_adapter_src_startofpacket                                                                                     : std_logic;                      -- width_adapter:out_startofpacket -> crosser_004:in_startofpacket
	signal width_adapter_src_data                                                                                              : std_logic_vector(90 downto 0);  -- width_adapter:out_data -> crosser_004:in_data
	signal width_adapter_src_ready                                                                                             : std_logic;                      -- crosser_004:in_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                                           : std_logic_vector(16 downto 0);  -- width_adapter:out_channel -> crosser_004:in_channel
	signal crosser_005_out_endofpacket                                                                                         : std_logic;                      -- crosser_005:out_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	signal crosser_005_out_valid                                                                                               : std_logic;                      -- crosser_005:out_valid -> cmd_xbar_mux_001:sink2_valid
	signal crosser_005_out_startofpacket                                                                                       : std_logic;                      -- crosser_005:out_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	signal crosser_005_out_data                                                                                                : std_logic_vector(90 downto 0);  -- crosser_005:out_data -> cmd_xbar_mux_001:sink2_data
	signal crosser_005_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_005:out_channel -> cmd_xbar_mux_001:sink2_channel
	signal crosser_005_out_ready                                                                                               : std_logic;                      -- cmd_xbar_mux_001:sink2_ready -> crosser_005:out_ready
	signal width_adapter_001_src_endofpacket                                                                                   : std_logic;                      -- width_adapter_001:out_endofpacket -> crosser_005:in_endofpacket
	signal width_adapter_001_src_valid                                                                                         : std_logic;                      -- width_adapter_001:out_valid -> crosser_005:in_valid
	signal width_adapter_001_src_startofpacket                                                                                 : std_logic;                      -- width_adapter_001:out_startofpacket -> crosser_005:in_startofpacket
	signal width_adapter_001_src_data                                                                                          : std_logic_vector(90 downto 0);  -- width_adapter_001:out_data -> crosser_005:in_data
	signal width_adapter_001_src_ready                                                                                         : std_logic;                      -- crosser_005:in_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                                       : std_logic_vector(16 downto 0);  -- width_adapter_001:out_channel -> crosser_005:in_channel
	signal crosser_006_out_endofpacket                                                                                         : std_logic;                      -- crosser_006:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal crosser_006_out_valid                                                                                               : std_logic;                      -- crosser_006:out_valid -> burst_adapter_001:sink0_valid
	signal crosser_006_out_startofpacket                                                                                       : std_logic;                      -- crosser_006:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal crosser_006_out_data                                                                                                : std_logic_vector(81 downto 0);  -- crosser_006:out_data -> burst_adapter_001:sink0_data
	signal crosser_006_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_006:out_channel -> burst_adapter_001:sink0_channel
	signal width_adapter_002_src_endofpacket                                                                                   : std_logic;                      -- width_adapter_002:out_endofpacket -> crosser_006:in_endofpacket
	signal width_adapter_002_src_valid                                                                                         : std_logic;                      -- width_adapter_002:out_valid -> crosser_006:in_valid
	signal width_adapter_002_src_startofpacket                                                                                 : std_logic;                      -- width_adapter_002:out_startofpacket -> crosser_006:in_startofpacket
	signal width_adapter_002_src_data                                                                                          : std_logic_vector(81 downto 0);  -- width_adapter_002:out_data -> crosser_006:in_data
	signal width_adapter_002_src_ready                                                                                         : std_logic;                      -- crosser_006:in_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                                       : std_logic_vector(16 downto 0);  -- width_adapter_002:out_channel -> crosser_006:in_channel
	signal crosser_007_out_endofpacket                                                                                         : std_logic;                      -- crosser_007:out_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal crosser_007_out_valid                                                                                               : std_logic;                      -- crosser_007:out_valid -> rsp_xbar_mux:sink1_valid
	signal crosser_007_out_startofpacket                                                                                       : std_logic;                      -- crosser_007:out_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal crosser_007_out_data                                                                                                : std_logic_vector(108 downto 0); -- crosser_007:out_data -> rsp_xbar_mux:sink1_data
	signal crosser_007_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_007:out_channel -> rsp_xbar_mux:sink1_channel
	signal crosser_007_out_ready                                                                                               : std_logic;                      -- rsp_xbar_mux:sink1_ready -> crosser_007:out_ready
	signal width_adapter_003_src_endofpacket                                                                                   : std_logic;                      -- width_adapter_003:out_endofpacket -> crosser_007:in_endofpacket
	signal width_adapter_003_src_valid                                                                                         : std_logic;                      -- width_adapter_003:out_valid -> crosser_007:in_valid
	signal width_adapter_003_src_startofpacket                                                                                 : std_logic;                      -- width_adapter_003:out_startofpacket -> crosser_007:in_startofpacket
	signal width_adapter_003_src_data                                                                                          : std_logic_vector(108 downto 0); -- width_adapter_003:out_data -> crosser_007:in_data
	signal width_adapter_003_src_ready                                                                                         : std_logic;                      -- crosser_007:in_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                                       : std_logic_vector(16 downto 0);  -- width_adapter_003:out_channel -> crosser_007:in_channel
	signal crosser_008_out_endofpacket                                                                                         : std_logic;                      -- crosser_008:out_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	signal crosser_008_out_valid                                                                                               : std_logic;                      -- crosser_008:out_valid -> rsp_xbar_mux_002:sink1_valid
	signal crosser_008_out_startofpacket                                                                                       : std_logic;                      -- crosser_008:out_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	signal crosser_008_out_data                                                                                                : std_logic_vector(108 downto 0); -- crosser_008:out_data -> rsp_xbar_mux_002:sink1_data
	signal crosser_008_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_008:out_channel -> rsp_xbar_mux_002:sink1_channel
	signal crosser_008_out_ready                                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink1_ready -> crosser_008:out_ready
	signal width_adapter_004_src_endofpacket                                                                                   : std_logic;                      -- width_adapter_004:out_endofpacket -> crosser_008:in_endofpacket
	signal width_adapter_004_src_valid                                                                                         : std_logic;                      -- width_adapter_004:out_valid -> crosser_008:in_valid
	signal width_adapter_004_src_startofpacket                                                                                 : std_logic;                      -- width_adapter_004:out_startofpacket -> crosser_008:in_startofpacket
	signal width_adapter_004_src_data                                                                                          : std_logic_vector(108 downto 0); -- width_adapter_004:out_data -> crosser_008:in_data
	signal width_adapter_004_src_ready                                                                                         : std_logic;                      -- crosser_008:in_ready -> width_adapter_004:out_ready
	signal width_adapter_004_src_channel                                                                                       : std_logic_vector(16 downto 0);  -- width_adapter_004:out_channel -> crosser_008:in_channel
	signal crosser_009_out_endofpacket                                                                                         : std_logic;                      -- crosser_009:out_endofpacket -> rsp_xbar_mux_002:sink7_endofpacket
	signal crosser_009_out_valid                                                                                               : std_logic;                      -- crosser_009:out_valid -> rsp_xbar_mux_002:sink7_valid
	signal crosser_009_out_startofpacket                                                                                       : std_logic;                      -- crosser_009:out_startofpacket -> rsp_xbar_mux_002:sink7_startofpacket
	signal crosser_009_out_data                                                                                                : std_logic_vector(108 downto 0); -- crosser_009:out_data -> rsp_xbar_mux_002:sink7_data
	signal crosser_009_out_channel                                                                                             : std_logic_vector(16 downto 0);  -- crosser_009:out_channel -> rsp_xbar_mux_002:sink7_channel
	signal crosser_009_out_ready                                                                                               : std_logic;                      -- rsp_xbar_mux_002:sink7_ready -> crosser_009:out_ready
	signal width_adapter_005_src_endofpacket                                                                                   : std_logic;                      -- width_adapter_005:out_endofpacket -> crosser_009:in_endofpacket
	signal width_adapter_005_src_valid                                                                                         : std_logic;                      -- width_adapter_005:out_valid -> crosser_009:in_valid
	signal width_adapter_005_src_startofpacket                                                                                 : std_logic;                      -- width_adapter_005:out_startofpacket -> crosser_009:in_startofpacket
	signal width_adapter_005_src_data                                                                                          : std_logic_vector(108 downto 0); -- width_adapter_005:out_data -> crosser_009:in_data
	signal width_adapter_005_src_ready                                                                                         : std_logic;                      -- crosser_009:in_ready -> width_adapter_005:out_ready
	signal width_adapter_005_src_channel                                                                                       : std_logic_vector(16 downto 0);  -- width_adapter_005:out_channel -> crosser_009:in_channel
	signal irq_mapper_receiver0_irq                                                                                            : std_logic;                      -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                                            : std_logic;                      -- sys_clk_timer:irq -> irq_mapper:receiver1_irq
	signal cpu_d_irq_irq                                                                                                       : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> cpu:d_irq
	signal reset_reset_n_ports_inv                                                                                             : std_logic;                      -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                                           : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart:av_read_n
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_write_ports_inv                                                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_anti_slave_0_write:inv -> sys_clk_timer:write_n
	signal red_led_pio_s1_translator_avalon_anti_slave_0_write_ports_inv                                                       : std_logic;                      -- red_led_pio_s1_translator_avalon_anti_slave_0_write:inv -> red_led_pio:write_n
	signal green_led_pio_s1_translator_avalon_anti_slave_0_write_ports_inv                                                     : std_logic;                      -- green_led_pio_s1_translator_avalon_anti_slave_0_write:inv -> green_led_pio:write_n
	signal control_out_s1_translator_avalon_anti_slave_0_write_ports_inv                                                       : std_logic;                      -- control_out_s1_translator_avalon_anti_slave_0_write:inv -> control_out:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                                            : std_logic;                      -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n]
	signal external_clocks_sys_clk_reset_reset_ports_inv                                                                       : std_logic;                      -- external_clocks_sys_clk_reset_reset:inv -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset_ports_inv                                                                        : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [FFT_in_0:reset_n, FFT_in_1:reset_n, FFT_in_2:reset_n, FFT_in_3:reset_n, control_in:reset_n, control_out:reset_n, green_led_pio:reset_n, red_led_pio:reset_n, rotary_in:reset_n, sys_clk_timer:reset_n, sysid:reset_n]

begin

	cpu : component nios2VGA_cpu
		port map (
			clk                                   => clk_clk,                                                          --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                         --                   reset_n.reset_n
			d_address                             => cpu_data_master_address,                                          --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                                       --                          .byteenable
			d_read                                => cpu_data_master_read,                                             --                          .read
			d_readdata                            => cpu_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => cpu_data_master_write,                                            --                          .write
			d_writedata                           => cpu_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                                   --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                                      --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                               --                          .waitrequest
			d_irq                                 => cpu_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                              -- custom_instruction_master.readra
		);

	jtag_uart : component nios2VGA_jtag_uart
		port map (
			clk            => clk_clk,                                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                   --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                    --               irq.irq
		);

	sys_clk_timer : component nios2VGA_sys_clk_timer
		port map (
			clk        => clk_clk,                                                         --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                    -- reset.reset_n
			address    => sys_clk_timer_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => sys_clk_timer_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                         --   irq.irq
		);

	sysid : component nios2VGA_sysid
		port map (
			clock    => clk_clk,                                                       --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,                  --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	red_led_pio : component nios2VGA_red_led_pio
		port map (
			clk        => clk_clk,                                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => red_led_pio_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => red_led_pio_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => red_led_pio_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => red_led_pio_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => red_led_pio_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => red_led_pio_external_connection_export                         -- external_connection.export
		);

	external_clocks : component nios2VGA_external_clocks
		port map (
			CLOCK_50    => clk_clk,                             --       clk_in_primary.clk
			reset       => rst_controller_001_reset_out_reset,  -- clk_in_primary_reset.reset
			sys_clk     => external_clocks_sys_clk_clk,         --              sys_clk.clk
			sys_reset_n => external_clocks_sys_clk_reset_reset, --        sys_clk_reset.reset_n
			SDRAM_CLK   => sdram_clock_clk,                     --            sdram_clk.clk
			VGA_CLK     => external_clocks_vga_clk_clk          --              vga_clk.clk
		);

	vga_dual_clock_fifo : component nios2VGA_VGA_Dual_Clock_FIFO
		port map (
			clk_stream_in            => external_clocks_sys_clk_clk,                               --         clock_stream_in.clk
			reset_stream_in          => rst_controller_002_reset_out_reset,                        --   clock_stream_in_reset.reset
			clk_stream_out           => external_clocks_vga_clk_clk,                               --        clock_stream_out.clk
			reset_stream_out         => rst_controller_003_reset_out_reset,                        --  clock_stream_out_reset.reset
			stream_in_ready          => alpha_blending_avalon_blended_source_ready,                --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => alpha_blending_avalon_blended_source_startofpacket,        --                        .startofpacket
			stream_in_endofpacket    => alpha_blending_avalon_blended_source_endofpacket,          --                        .endofpacket
			stream_in_valid          => alpha_blending_avalon_blended_source_valid,                --                        .valid
			stream_in_data           => alpha_blending_avalon_blended_source_data,                 --                        .data
			stream_out_ready         => vga_dual_clock_fifo_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => vga_dual_clock_fifo_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => vga_dual_clock_fifo_avalon_dc_buffer_source_data           --                        .data
		);

	alpha_blending : component nios2VGA_Alpha_Blending
		port map (
			clk                      => external_clocks_sys_clk_clk,                           --            clock_reset.clk
			reset                    => rst_controller_002_reset_out_reset,                    --      clock_reset_reset.reset
			foreground_data          => vga_character_buffer_avalon_char_source_data,          -- avalon_foreground_sink.data
			foreground_startofpacket => vga_character_buffer_avalon_char_source_startofpacket, --                       .startofpacket
			foreground_endofpacket   => vga_character_buffer_avalon_char_source_endofpacket,   --                       .endofpacket
			foreground_valid         => vga_character_buffer_avalon_char_source_valid,         --                       .valid
			foreground_ready         => vga_character_buffer_avalon_char_source_ready,         --                       .ready
			background_data          => vga_scaler_avalon_scaler_source_data,                  -- avalon_background_sink.data
			background_startofpacket => vga_scaler_avalon_scaler_source_startofpacket,         --                       .startofpacket
			background_endofpacket   => vga_scaler_avalon_scaler_source_endofpacket,           --                       .endofpacket
			background_valid         => vga_scaler_avalon_scaler_source_valid,                 --                       .valid
			background_ready         => vga_scaler_avalon_scaler_source_ready,                 --                       .ready
			output_ready             => alpha_blending_avalon_blended_source_ready,            --  avalon_blended_source.ready
			output_data              => alpha_blending_avalon_blended_source_data,             --                       .data
			output_startofpacket     => alpha_blending_avalon_blended_source_startofpacket,    --                       .startofpacket
			output_endofpacket       => alpha_blending_avalon_blended_source_endofpacket,      --                       .endofpacket
			output_valid             => alpha_blending_avalon_blended_source_valid             --                       .valid
		);

	vga_controller : component nios2VGA_VGA_Controller
		port map (
			clk           => external_clocks_vga_clk_clk,                               --        clock_reset.clk
			reset         => rst_controller_003_reset_out_reset,                        --  clock_reset_reset.reset
			data          => vga_dual_clock_fifo_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => vga_dual_clock_fifo_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => vga_dual_clock_fifo_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_controller_external_CLK,                               -- external_interface.export
			VGA_HS        => vga_controller_external_HS,                                --                   .export
			VGA_VS        => vga_controller_external_VS,                                --                   .export
			VGA_BLANK     => vga_controller_external_BLANK,                             --                   .export
			VGA_SYNC      => vga_controller_external_SYNC,                              --                   .export
			VGA_R         => vga_controller_external_R,                                 --                   .export
			VGA_G         => vga_controller_external_G,                                 --                   .export
			VGA_B         => vga_controller_external_B                                  --                   .export
		);

	vga_character_buffer : component nios2VGA_VGA_Character_buffer
		port map (
			clk                  => external_clocks_sys_clk_clk,                                                                --               clock_reset.clk
			reset                => rst_controller_002_reset_out_reset,                                                         --         clock_reset_reset.reset
			ctrl_address         => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address(0),   -- avalon_char_control_slave.address
			ctrl_byteenable      => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable,   --                          .byteenable
			ctrl_chipselect      => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect,   --                          .chipselect
			ctrl_read            => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read,         --                          .read
			ctrl_write           => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write,        --                          .write
			ctrl_writedata       => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata,    --                          .writedata
			ctrl_readdata        => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata,     --                          .readdata
			buf_byteenable       => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable(0), --  avalon_char_buffer_slave.byteenable
			buf_chipselect       => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect,    --                          .chipselect
			buf_read             => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read,          --                          .read
			buf_write            => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write,         --                          .write
			buf_writedata        => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata,     --                          .writedata
			buf_readdata         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata,      --                          .readdata
			buf_waitrequest      => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest,   --                          .waitrequest
			buf_address          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address,       --                          .address
			stream_ready         => vga_character_buffer_avalon_char_source_ready,                                              --        avalon_char_source.ready
			stream_startofpacket => vga_character_buffer_avalon_char_source_startofpacket,                                      --                          .startofpacket
			stream_endofpacket   => vga_character_buffer_avalon_char_source_endofpacket,                                        --                          .endofpacket
			stream_valid         => vga_character_buffer_avalon_char_source_valid,                                              --                          .valid
			stream_data          => vga_character_buffer_avalon_char_source_data                                                --                          .data
		);

	vga_scaler : component nios2VGA_VGA_Scaler
		port map (
			clk                      => external_clocks_sys_clk_clk,                             --          clock_reset.clk
			reset                    => rst_controller_002_reset_out_reset,                      --    clock_reset_reset.reset
			stream_in_startofpacket  => vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => vga_pixel_rgb_resampler_avalon_rgb_source_valid,         --                     .valid
			stream_in_ready          => vga_pixel_rgb_resampler_avalon_rgb_source_ready,         --                     .ready
			stream_in_data           => vga_pixel_rgb_resampler_avalon_rgb_source_data,          --                     .data
			stream_out_ready         => vga_scaler_avalon_scaler_source_ready,                   -- avalon_scaler_source.ready
			stream_out_startofpacket => vga_scaler_avalon_scaler_source_startofpacket,           --                     .startofpacket
			stream_out_endofpacket   => vga_scaler_avalon_scaler_source_endofpacket,             --                     .endofpacket
			stream_out_valid         => vga_scaler_avalon_scaler_source_valid,                   --                     .valid
			stream_out_data          => vga_scaler_avalon_scaler_source_data                     --                     .data
		);

	vga_pixel_rgb_resampler : component nios2VGA_VGA_pixel_RGB_Resampler
		port map (
			clk                      => external_clocks_sys_clk_clk,                             --       clock_reset.clk
			reset                    => rst_controller_002_reset_out_reset,                      -- clock_reset_reset.reset
			stream_in_startofpacket  => vga_pixel_buffer_avalon_pixel_source_startofpacket,      --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => vga_pixel_buffer_avalon_pixel_source_endofpacket,        --                  .endofpacket
			stream_in_valid          => vga_pixel_buffer_avalon_pixel_source_valid,              --                  .valid
			stream_in_ready          => vga_pixel_buffer_avalon_pixel_source_ready,              --                  .ready
			stream_in_data           => vga_pixel_buffer_avalon_pixel_source_data,               --                  .data
			stream_out_ready         => vga_pixel_rgb_resampler_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => vga_pixel_rgb_resampler_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => vga_pixel_rgb_resampler_avalon_rgb_source_data           --                  .data
		);

	vga_pixel_buffer : component nios2VGA_VGA_Pixel_Buffer
		port map (
			clk                  => external_clocks_sys_clk_clk,                                                     --             clock_reset.clk
			reset                => rst_controller_002_reset_out_reset,                                              --       clock_reset_reset.reset
			master_readdatavalid => vga_pixel_buffer_avalon_pixel_dma_master_readdatavalid,                          -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => vga_pixel_buffer_avalon_pixel_dma_master_waitrequest,                            --                        .waitrequest
			master_address       => vga_pixel_buffer_avalon_pixel_dma_master_address,                                --                        .address
			master_arbiterlock   => vga_pixel_buffer_avalon_pixel_dma_master_lock,                                   --                        .lock
			master_read          => vga_pixel_buffer_avalon_pixel_dma_master_read,                                   --                        .read
			master_readdata      => vga_pixel_buffer_avalon_pixel_dma_master_readdata,                               --                        .readdata
			slave_address        => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_address,    --    avalon_control_slave.address
			slave_byteenable     => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_byteenable, --                        .byteenable
			slave_read           => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_read,       --                        .read
			slave_write          => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_write,      --                        .write
			slave_writedata      => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_writedata,  --                        .writedata
			slave_readdata       => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_readdata,   --                        .readdata
			stream_ready         => vga_pixel_buffer_avalon_pixel_source_ready,                                      --     avalon_pixel_source.ready
			stream_startofpacket => vga_pixel_buffer_avalon_pixel_source_startofpacket,                              --                        .startofpacket
			stream_endofpacket   => vga_pixel_buffer_avalon_pixel_source_endofpacket,                                --                        .endofpacket
			stream_valid         => vga_pixel_buffer_avalon_pixel_source_valid,                                      --                        .valid
			stream_data          => vga_pixel_buffer_avalon_pixel_source_data                                        --                        .data
		);

	sram : component nios2VGA_SRAM
		port map (
			clk           => external_clocks_sys_clk_clk,                                         --        clock_reset.clk
			reset         => rst_controller_002_reset_out_reset,                                  --  clock_reset_reset.reset
			SRAM_DQ       => sram_external_interface_DQ,                                          -- external_interface.export
			SRAM_ADDR     => sram_external_interface_ADDR,                                        --                   .export
			SRAM_LB_N     => sram_external_interface_LB_N,                                        --                   .export
			SRAM_UB_N     => sram_external_interface_UB_N,                                        --                   .export
			SRAM_CE_N     => sram_external_interface_CE_N,                                        --                   .export
			SRAM_OE_N     => sram_external_interface_OE_N,                                        --                   .export
			SRAM_WE_N     => sram_external_interface_WE_N,                                        --                   .export
			address       => sram_avalon_sram_slave_translator_avalon_anti_slave_0_address,       --  avalon_sram_slave.address
			byteenable    => sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,    --                   .byteenable
			read          => sram_avalon_sram_slave_translator_avalon_anti_slave_0_read,          --                   .read
			write         => sram_avalon_sram_slave_translator_avalon_anti_slave_0_write,         --                   .write
			writedata     => sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,     --                   .writedata
			readdata      => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,      --                   .readdata
			readdatavalid => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid  --                   .readdatavalid
		);

	green_led_pio : component nios2VGA_green_led_pio
		port map (
			clk        => clk_clk,                                                         --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => green_led_pio_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => green_led_pio_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => green_led_pio_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => green_led_pio_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => green_led_pio_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => green_led_pio_external_connection_export                         -- external_connection.export
		);

	control_in : component nios2VGA_control_in
		port map (
			clk      => clk_clk,                                               --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,          --               reset.reset_n
			address  => control_in_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => control_in_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => nios_cntrl_in_export                                   -- external_connection.export
		);

	control_out : component nios2VGA_control_out
		port map (
			clk        => clk_clk,                                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => control_out_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => control_out_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => control_out_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => control_out_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => control_out_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => nios_cntrl_out_export                                          -- external_connection.export
		);

	fft_in_0 : component nios2VGA_FFT_in_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,        --               reset.reset_n
			address  => fft_in_0_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => fft_in_0_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => fft_in_0_export                                      -- external_connection.export
		);

	fft_in_1 : component nios2VGA_FFT_in_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,        --               reset.reset_n
			address  => fft_in_1_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => fft_in_1_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => fft_in_1_export                                      -- external_connection.export
		);

	fft_in_2 : component nios2VGA_FFT_in_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,        --               reset.reset_n
			address  => fft_in_2_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => fft_in_2_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => fft_in_2_export                                      -- external_connection.export
		);

	fft_in_3 : component nios2VGA_FFT_in_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,        --               reset.reset_n
			address  => fft_in_3_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => fft_in_3_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => fft_in_3_export                                      -- external_connection.export
		);

	rotary_in : component nios2VGA_control_in
		port map (
			clk      => clk_clk,                                              --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address  => rotary_in_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => rotary_in_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => rotary_in_export                                      -- external_connection.export
		);

	cpu_instruction_master_translator : component nios2vga_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 20,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                   --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                       --               (terminated)
			av_byteenable            => "1111",                                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_readdatavalid         => open,                                                                      --               (terminated)
			av_write                 => '0',                                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			av_debugaccess           => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	vga_pixel_buffer_avalon_pixel_dma_master_translator : component nios2vga_vga_pixel_buffer_avalon_pixel_dma_master_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 16,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 2,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 2,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 2,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                                 --                       clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                          --                     reset.reset
			uav_address              => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => vga_pixel_buffer_avalon_pixel_dma_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => vga_pixel_buffer_avalon_pixel_dma_master_waitrequest,                                        --                          .waitrequest
			av_read                  => vga_pixel_buffer_avalon_pixel_dma_master_read,                                               --                          .read
			av_readdata              => vga_pixel_buffer_avalon_pixel_dma_master_readdata,                                           --                          .readdata
			av_readdatavalid         => vga_pixel_buffer_avalon_pixel_dma_master_readdatavalid,                                      --                          .readdatavalid
			av_lock                  => vga_pixel_buffer_avalon_pixel_dma_master_lock,                                               --                          .lock
			av_burstcount            => "1",                                                                                         --               (terminated)
			av_byteenable            => "11",                                                                                        --               (terminated)
			av_beginbursttransfer    => '0',                                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                                         --               (terminated)
			av_chipselect            => '0',                                                                                         --               (terminated)
			av_write                 => '0',                                                                                         --               (terminated)
			av_writedata             => "0000000000000000",                                                                          --               (terminated)
			av_debugaccess           => '0',                                                                                         --               (terminated)
			uav_clken                => open,                                                                                        --               (terminated)
			av_clken                 => '1',                                                                                         --               (terminated)
			uav_response             => "00",                                                                                        --               (terminated)
			av_response              => open,                                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                                         --               (terminated)
		);

	cpu_data_master_translator : component nios2vga_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 20,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clk_clk,                                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_data_master_read,                                               --                          .read
			av_readdata              => cpu_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_data_master_write,                                              --                          .write
			av_writedata             => cpu_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_readdatavalid         => open,                                                               --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	cpu_jtag_debug_module_translator : component nios2vga_cpu_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_chipselect            => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	sram_avalon_sram_slave_translator : component nios2vga_sram_avalon_sram_slave_translator
		generic map (
			AV_ADDRESS_W                   => 18,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                       --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                --                    reset.reset
			uav_address              => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sram_avalon_sram_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sram_avalon_sram_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sram_avalon_sram_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_chipselect            => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator : component nios2vga_jtag_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	sys_clk_timer_s1_translator : component nios2vga_sys_clk_timer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                     --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                          --                    reset.reset
			uav_address              => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sys_clk_timer_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sys_clk_timer_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	sysid_control_slave_translator : component nios2vga_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                             --                    reset.reset
			uav_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                           --              (terminated)
			av_read                  => open,                                                                           --              (terminated)
			av_writedata             => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	red_led_pio_s1_translator : component nios2vga_red_led_pio_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                   --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                        --                    reset.reset
			uav_address              => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => red_led_pio_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => red_led_pio_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => red_led_pio_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => red_led_pio_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => red_led_pio_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                      --              (terminated)
			av_begintransfer         => open,                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                      --              (terminated)
			av_burstcount            => open,                                                                      --              (terminated)
			av_byteenable            => open,                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                      --              (terminated)
			av_lock                  => open,                                                                      --              (terminated)
			av_clken                 => open,                                                                      --              (terminated)
			uav_clken                => '0',                                                                       --              (terminated)
			av_debugaccess           => open,                                                                      --              (terminated)
			av_outputenable          => open,                                                                      --              (terminated)
			uav_response             => open,                                                                      --              (terminated)
			av_response              => "00",                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                        --              (terminated)
		);

	vga_character_buffer_avalon_char_control_slave_translator : component nios2vga_vga_character_buffer_avalon_char_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                                               --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                                        --                    reset.reset
			uav_address              => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                                      --              (terminated)
			av_lock                  => open,                                                                                                      --              (terminated)
			av_clken                 => open,                                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                                      --              (terminated)
			uav_response             => open,                                                                                                      --              (terminated)
			av_response              => "00",                                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                                        --              (terminated)
		);

	vga_character_buffer_avalon_char_buffer_slave_translator : component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator
		generic map (
			AV_ADDRESS_W                   => 13,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 8,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 1,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 1,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 1,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                                              --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                                       --                    reset.reset
			uav_address              => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                                                     --              (terminated)
			av_burstcount            => open,                                                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                                                     --              (terminated)
			av_lock                  => open,                                                                                                     --              (terminated)
			av_clken                 => open,                                                                                                     --              (terminated)
			uav_clken                => '0',                                                                                                      --              (terminated)
			av_debugaccess           => open,                                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                                     --              (terminated)
			uav_response             => open,                                                                                                     --              (terminated)
			av_response              => "00",                                                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                                                       --              (terminated)
		);

	vga_pixel_buffer_avalon_control_slave_translator : component nios2vga_vga_pixel_buffer_avalon_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                                      --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                               --                    reset.reset
			uav_address              => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_begintransfer         => open,                                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                                             --              (terminated)
			av_burstcount            => open,                                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                                             --              (terminated)
			av_lock                  => open,                                                                                             --              (terminated)
			av_chipselect            => open,                                                                                             --              (terminated)
			av_clken                 => open,                                                                                             --              (terminated)
			uav_clken                => '0',                                                                                              --              (terminated)
			av_debugaccess           => open,                                                                                             --              (terminated)
			av_outputenable          => open,                                                                                             --              (terminated)
			uav_response             => open,                                                                                             --              (terminated)
			av_response              => "00",                                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                                               --              (terminated)
		);

	green_led_pio_s1_translator : component nios2vga_red_led_pio_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                     --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                          --                    reset.reset
			uav_address              => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => green_led_pio_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => green_led_pio_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => green_led_pio_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => green_led_pio_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => green_led_pio_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	control_in_s1_translator : component nios2vga_control_in_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                       --                    reset.reset
			uav_address              => control_in_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => control_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => control_in_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => control_in_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => control_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => control_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => control_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => control_in_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => control_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => control_in_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => control_in_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                     --              (terminated)
			av_read                  => open,                                                                     --              (terminated)
			av_writedata             => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_chipselect            => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	control_out_s1_translator : component nios2vga_red_led_pio_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                   --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                        --                    reset.reset
			uav_address              => control_out_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => control_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => control_out_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => control_out_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => control_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => control_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => control_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => control_out_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => control_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => control_out_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => control_out_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => control_out_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => control_out_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => control_out_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                      --              (terminated)
			av_begintransfer         => open,                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                      --              (terminated)
			av_burstcount            => open,                                                                      --              (terminated)
			av_byteenable            => open,                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                      --              (terminated)
			av_lock                  => open,                                                                      --              (terminated)
			av_clken                 => open,                                                                      --              (terminated)
			uav_clken                => '0',                                                                       --              (terminated)
			av_debugaccess           => open,                                                                      --              (terminated)
			av_outputenable          => open,                                                                      --              (terminated)
			uav_response             => open,                                                                      --              (terminated)
			av_response              => "00",                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                        --              (terminated)
		);

	fft_in_0_s1_translator : component nios2vga_control_in_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                     --                    reset.reset
			uav_address              => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => fft_in_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => fft_in_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                   --              (terminated)
			av_read                  => open,                                                                   --              (terminated)
			av_writedata             => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_chipselect            => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	fft_in_1_s1_translator : component nios2vga_control_in_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                     --                    reset.reset
			uav_address              => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => fft_in_1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => fft_in_1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                   --              (terminated)
			av_read                  => open,                                                                   --              (terminated)
			av_writedata             => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_chipselect            => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	fft_in_2_s1_translator : component nios2vga_control_in_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                     --                    reset.reset
			uav_address              => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => fft_in_2_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => fft_in_2_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                   --              (terminated)
			av_read                  => open,                                                                   --              (terminated)
			av_writedata             => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_chipselect            => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	fft_in_3_s1_translator : component nios2vga_control_in_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                     --                    reset.reset
			uav_address              => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => fft_in_3_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => fft_in_3_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                   --              (terminated)
			av_read                  => open,                                                                   --              (terminated)
			av_writedata             => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_chipselect            => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	rotary_in_s1_translator : component nios2vga_control_in_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                 --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                      --                    reset.reset
			uav_address              => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => rotary_in_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => rotary_in_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                    --              (terminated)
			av_read                  => open,                                                                    --              (terminated)
			av_writedata             => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_chipselect            => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	cpu_instruction_master_translator_avalon_universal_master_0_agent : component nios2vga_cpu_instruction_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_BEGIN_BURST           => 87,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			PKT_BURST_TYPE_H          => 84,
			PKT_BURST_TYPE_L          => 83,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_THREAD_ID_H           => 99,
			PKT_THREAD_ID_L           => 99,
			PKT_CACHE_H               => 106,
			PKT_CACHE_L               => 103,
			PKT_DATA_SIDEBAND_H       => 86,
			PKT_DATA_SIDEBAND_L       => 86,
			PKT_QOS_H                 => 88,
			PKT_QOS_L                 => 88,
			PKT_ADDR_SIDEBAND_H       => 85,
			PKT_ADDR_SIDEBAND_L       => 85,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			ST_DATA_W                 => 109,
			ST_CHANNEL_W              => 17,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 2,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                            --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                             --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                              --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                           --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                     --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                       --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                             --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent : component nios2vga_vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 84,
			PKT_PROTECTION_L          => 82,
			PKT_BEGIN_BURST           => 69,
			PKT_BURSTWRAP_H           => 61,
			PKT_BURSTWRAP_L           => 59,
			PKT_BURST_SIZE_H          => 64,
			PKT_BURST_SIZE_L          => 62,
			PKT_BURST_TYPE_H          => 66,
			PKT_BURST_TYPE_L          => 65,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_TRANS_EXCLUSIVE       => 55,
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 71,
			PKT_DEST_ID_H             => 80,
			PKT_DEST_ID_L             => 76,
			PKT_THREAD_ID_H           => 81,
			PKT_THREAD_ID_L           => 81,
			PKT_CACHE_H               => 88,
			PKT_CACHE_L               => 85,
			PKT_DATA_SIDEBAND_H       => 68,
			PKT_DATA_SIDEBAND_L       => 68,
			PKT_QOS_H                 => 70,
			PKT_QOS_L                 => 70,
			PKT_ADDR_SIDEBAND_H       => 67,
			PKT_ADDR_SIDEBAND_L       => 67,
			PKT_RESPONSE_STATUS_H     => 90,
			PKT_RESPONSE_STATUS_L     => 89,
			ST_DATA_W                 => 91,
			ST_CHANNEL_W              => 17,
			AV_BURSTCOUNT_W           => 2,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                          --       clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                                   -- clk_reset.reset
			av_address              => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_001_src1_valid,                                                                        --        rp.valid
			rp_data                 => rsp_xbar_demux_001_src1_data,                                                                         --          .data
			rp_channel              => rsp_xbar_demux_001_src1_channel,                                                                      --          .channel
			rp_startofpacket        => rsp_xbar_demux_001_src1_startofpacket,                                                                --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_001_src1_endofpacket,                                                                  --          .endofpacket
			rp_ready                => rsp_xbar_demux_001_src1_ready,                                                                        --          .ready
			av_response             => open,                                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                                  -- (terminated)
		);

	cpu_data_master_translator_avalon_universal_master_0_agent : component nios2vga_cpu_instruction_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_BEGIN_BURST           => 87,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			PKT_BURST_TYPE_H          => 84,
			PKT_BURST_TYPE_L          => 83,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_THREAD_ID_H           => 99,
			PKT_THREAD_ID_L           => 99,
			PKT_CACHE_H               => 106,
			PKT_CACHE_L               => 103,
			PKT_DATA_SIDEBAND_H       => 86,
			PKT_DATA_SIDEBAND_L       => 86,
			PKT_QOS_H                 => 88,
			PKT_QOS_L                 => 88,
			PKT_ADDR_SIDEBAND_H       => 85,
			PKT_ADDR_SIDEBAND_L       => 85,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			ST_DATA_W                 => 109,
			ST_CHANNEL_W              => 17,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_002_src_valid,                                                  --        rp.valid
			rp_data                 => rsp_xbar_mux_002_src_data,                                                   --          .data
			rp_channel              => rsp_xbar_mux_002_src_channel,                                                --          .channel
			rp_startofpacket        => rsp_xbar_mux_002_src_startofpacket,                                          --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_002_src_endofpacket,                                            --          .endofpacket
			rp_ready                => rsp_xbar_mux_002_src_ready,                                                  --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                     --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                   --                .channel
			rf_sink_ready           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                 -- (terminated)
			csr_read          => '0',                                                                                  -- (terminated)
			csr_write         => '0',                                                                                  -- (terminated)
			csr_readdata      => open,                                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                   -- (terminated)
			almost_full_data  => open,                                                                                 -- (terminated)
			almost_empty_data => open,                                                                                 -- (terminated)
			in_startofpacket  => '0',                                                                                  -- (terminated)
			in_endofpacket    => '0',                                                                                  -- (terminated)
			out_startofpacket => open,                                                                                 -- (terminated)
			out_endofpacket   => open,                                                                                 -- (terminated)
			in_empty          => '0',                                                                                  -- (terminated)
			out_empty         => open,                                                                                 -- (terminated)
			in_error          => '0',                                                                                  -- (terminated)
			out_error         => open,                                                                                 -- (terminated)
			in_channel        => '0',                                                                                  -- (terminated)
			out_channel       => open                                                                                  -- (terminated)
		);

	sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent : component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 69,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 71,
			PKT_DEST_ID_H             => 80,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 61,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 84,
			PKT_PROTECTION_L          => 82,
			PKT_RESPONSE_STATUS_H     => 90,
			PKT_RESPONSE_STATUS_L     => 89,
			PKT_BURST_SIZE_H          => 64,
			PKT_BURST_SIZE_L          => 62,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 91,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                 --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                 --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                 --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                  --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                         --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                           --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                               --                .channel
			rf_sink_ready           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 92,
			FIFO_DEPTH          => 3,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                 --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 3,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                           --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_startofpacket  => '0',                                                                                   -- (terminated)
			in_endofpacket    => '0',                                                                                   -- (terminated)
			out_startofpacket => open,                                                                                  -- (terminated)
			out_endofpacket   => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src2_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src2_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_demux_002_src2_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src2_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src2_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src2_channel,                                                                  --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_startofpacket  => '0',                                                                                        -- (terminated)
			in_endofpacket    => '0',                                                                                        -- (terminated)
			out_startofpacket => open,                                                                                       -- (terminated)
			out_endofpacket   => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	sys_clk_timer_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                               --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src3_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src3_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_demux_002_src3_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src3_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src3_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src3_channel,                                                       --                .channel
			rf_sink_ready           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                               --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_startofpacket  => '0',                                                                             -- (terminated)
			in_endofpacket    => '0',                                                                             -- (terminated)
			out_startofpacket => open,                                                                            -- (terminated)
			out_endofpacket   => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                       --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src4_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src4_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_002_src4_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src4_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src4_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src4_channel,                                                          --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_startofpacket  => '0',                                                                                -- (terminated)
			in_endofpacket    => '0',                                                                                -- (terminated)
			out_startofpacket => open,                                                                               -- (terminated)
			out_endofpacket   => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	red_led_pio_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                             --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src5_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src5_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_demux_002_src5_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src5_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src5_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src5_channel,                                                     --                .channel
			rf_sink_ready           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                  --     (terminated)
		);

	red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                             --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                -- (terminated)
			csr_read          => '0',                                                                                 -- (terminated)
			csr_write         => '0',                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                  -- (terminated)
			almost_full_data  => open,                                                                                -- (terminated)
			almost_empty_data => open,                                                                                -- (terminated)
			in_empty          => '0',                                                                                 -- (terminated)
			out_empty         => open,                                                                                -- (terminated)
			in_error          => '0',                                                                                 -- (terminated)
			out_error         => open,                                                                                -- (terminated)
			in_channel        => '0',                                                                                 -- (terminated)
			out_channel       => open                                                                                 -- (terminated)
		);

	red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                       --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			in_data           => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_startofpacket  => '0',                                                                           -- (terminated)
			in_endofpacket    => '0',                                                                           -- (terminated)
			out_startofpacket => open,                                                                          -- (terminated)
			out_endofpacket   => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                                         --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                                                  --       clk_reset.reset
			m0_address              => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => crosser_out_ready,                                                                                                   --              cp.ready
			cp_valid                => crosser_out_valid,                                                                                                   --                .valid
			cp_data                 => crosser_out_data,                                                                                                    --                .data
			cp_startofpacket        => crosser_out_startofpacket,                                                                                           --                .startofpacket
			cp_endofpacket          => crosser_out_endofpacket,                                                                                             --                .endofpacket
			cp_channel              => crosser_out_channel,                                                                                                 --                .channel
			rf_sink_ready           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                                  --     (terminated)
		);

	vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                                         --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                                                  -- clk_reset.reset
			in_data           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                                -- (terminated)
			in_error          => '0',                                                                                                                 -- (terminated)
			out_error         => open,                                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                                 -- (terminated)
			out_channel       => open                                                                                                                 -- (terminated)
		);

	vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                                   --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                                            -- clk_reset.reset
			in_data           => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                                          -- (terminated)
			csr_read          => '0',                                                                                                           -- (terminated)
			csr_write         => '0',                                                                                                           -- (terminated)
			csr_readdata      => open,                                                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                            -- (terminated)
			almost_full_data  => open,                                                                                                          -- (terminated)
			almost_empty_data => open,                                                                                                          -- (terminated)
			in_startofpacket  => '0',                                                                                                           -- (terminated)
			in_endofpacket    => '0',                                                                                                           -- (terminated)
			out_startofpacket => open,                                                                                                          -- (terminated)
			out_endofpacket   => open,                                                                                                          -- (terminated)
			in_empty          => '0',                                                                                                           -- (terminated)
			out_empty         => open,                                                                                                          -- (terminated)
			in_error          => '0',                                                                                                           -- (terminated)
			out_error         => open,                                                                                                          -- (terminated)
			in_channel        => '0',                                                                                                           -- (terminated)
			out_channel       => open                                                                                                           -- (terminated)
		);

	vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent : component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 7,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 60,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_POSTED          => 42,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			PKT_TRANS_LOCK            => 45,
			PKT_SRC_ID_H              => 66,
			PKT_SRC_ID_L              => 62,
			PKT_DEST_ID_H             => 71,
			PKT_DEST_ID_L             => 67,
			PKT_BURSTWRAP_H           => 52,
			PKT_BURSTWRAP_L           => 50,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_PROTECTION_H          => 75,
			PKT_PROTECTION_L          => 73,
			PKT_RESPONSE_STATUS_H     => 81,
			PKT_RESPONSE_STATUS_L     => 80,
			PKT_BURST_SIZE_H          => 55,
			PKT_BURST_SIZE_L          => 53,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 82,
			AVS_BURSTCOUNT_W          => 1,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                                        --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                                                 --       clk_reset.reset
			m0_address              => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                                                    --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                                                    --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                                                     --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                                                            --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                                                              --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                                                  --                .channel
			rf_sink_ready           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                                 --     (terminated)
		);

	vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 83,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                                        --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                                                 -- clk_reset.reset
			in_data           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                               -- (terminated)
			csr_read          => '0',                                                                                                                -- (terminated)
			csr_write         => '0',                                                                                                                -- (terminated)
			csr_readdata      => open,                                                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                                 -- (terminated)
			almost_full_data  => open,                                                                                                               -- (terminated)
			almost_empty_data => open,                                                                                                               -- (terminated)
			in_empty          => '0',                                                                                                                -- (terminated)
			out_empty         => open,                                                                                                               -- (terminated)
			in_error          => '0',                                                                                                                -- (terminated)
			out_error         => open,                                                                                                               -- (terminated)
			in_channel        => '0',                                                                                                                -- (terminated)
			out_channel       => open                                                                                                                -- (terminated)
		);

	vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 10,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                                           -- clk_reset.reset
			in_data           => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                                         -- (terminated)
			csr_read          => '0',                                                                                                          -- (terminated)
			csr_write         => '0',                                                                                                          -- (terminated)
			csr_readdata      => open,                                                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                           -- (terminated)
			almost_full_data  => open,                                                                                                         -- (terminated)
			almost_empty_data => open,                                                                                                         -- (terminated)
			in_startofpacket  => '0',                                                                                                          -- (terminated)
			in_endofpacket    => '0',                                                                                                          -- (terminated)
			out_startofpacket => open,                                                                                                         -- (terminated)
			out_endofpacket   => open,                                                                                                         -- (terminated)
			in_empty          => '0',                                                                                                          -- (terminated)
			out_empty         => open,                                                                                                         -- (terminated)
			in_error          => '0',                                                                                                          -- (terminated)
			out_error         => open,                                                                                                         -- (terminated)
			in_channel        => '0',                                                                                                          -- (terminated)
			out_channel       => open                                                                                                          -- (terminated)
		);

	vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                                --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                                         --       clk_reset.reset
			m0_address              => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => crosser_001_out_ready,                                                                                      --              cp.ready
			cp_valid                => crosser_001_out_valid,                                                                                      --                .valid
			cp_data                 => crosser_001_out_data,                                                                                       --                .data
			cp_startofpacket        => crosser_001_out_startofpacket,                                                                              --                .startofpacket
			cp_endofpacket          => crosser_001_out_endofpacket,                                                                                --                .endofpacket
			cp_channel              => crosser_001_out_channel,                                                                                    --                .channel
			rf_sink_ready           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                         --     (terminated)
		);

	vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                                --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                                         -- clk_reset.reset
			in_data           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                       -- (terminated)
			csr_read          => '0',                                                                                                        -- (terminated)
			csr_write         => '0',                                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                         -- (terminated)
			almost_full_data  => open,                                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                                       -- (terminated)
			in_empty          => '0',                                                                                                        -- (terminated)
			out_empty         => open,                                                                                                       -- (terminated)
			in_error          => '0',                                                                                                        -- (terminated)
			out_error         => open,                                                                                                       -- (terminated)
			in_channel        => '0',                                                                                                        -- (terminated)
			out_channel       => open                                                                                                        -- (terminated)
		);

	vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                                 -- (terminated)
			csr_read          => '0',                                                                                                  -- (terminated)
			csr_write         => '0',                                                                                                  -- (terminated)
			csr_readdata      => open,                                                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                   -- (terminated)
			almost_full_data  => open,                                                                                                 -- (terminated)
			almost_empty_data => open,                                                                                                 -- (terminated)
			in_startofpacket  => '0',                                                                                                  -- (terminated)
			in_endofpacket    => '0',                                                                                                  -- (terminated)
			out_startofpacket => open,                                                                                                 -- (terminated)
			out_endofpacket   => open,                                                                                                 -- (terminated)
			in_empty          => '0',                                                                                                  -- (terminated)
			out_empty         => open,                                                                                                 -- (terminated)
			in_error          => '0',                                                                                                  -- (terminated)
			out_error         => open,                                                                                                 -- (terminated)
			in_channel        => '0',                                                                                                  -- (terminated)
			out_channel       => open                                                                                                  -- (terminated)
		);

	green_led_pio_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                               --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src9_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src9_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_demux_002_src9_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src9_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src9_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src9_channel,                                                       --                .channel
			rf_sink_ready           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                               --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_startofpacket  => '0',                                                                             -- (terminated)
			in_endofpacket    => '0',                                                                             -- (terminated)
			out_startofpacket => open,                                                                            -- (terminated)
			out_endofpacket   => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	control_in_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                            --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => control_in_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => control_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => control_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => control_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => control_in_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => control_in_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => control_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => control_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => control_in_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => control_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => control_in_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => control_in_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => control_in_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => control_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src10_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src10_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_002_src10_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src10_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src10_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src10_channel,                                                   --                .channel
			rf_sink_ready           => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                           -- clk_reset.reset
			in_data           => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                         -- (terminated)
			csr_read          => '0',                                                                          -- (terminated)
			csr_write         => '0',                                                                          -- (terminated)
			csr_readdata      => open,                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                           -- (terminated)
			almost_full_data  => open,                                                                         -- (terminated)
			almost_empty_data => open,                                                                         -- (terminated)
			in_startofpacket  => '0',                                                                          -- (terminated)
			in_endofpacket    => '0',                                                                          -- (terminated)
			out_startofpacket => open,                                                                         -- (terminated)
			out_endofpacket   => open,                                                                         -- (terminated)
			in_empty          => '0',                                                                          -- (terminated)
			out_empty         => open,                                                                         -- (terminated)
			in_error          => '0',                                                                          -- (terminated)
			out_error         => open,                                                                         -- (terminated)
			in_channel        => '0',                                                                          -- (terminated)
			out_channel       => open                                                                          -- (terminated)
		);

	control_out_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                             --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => control_out_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => control_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => control_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => control_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => control_out_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => control_out_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => control_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => control_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => control_out_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => control_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => control_out_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => control_out_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => control_out_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => control_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src11_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src11_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_demux_002_src11_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src11_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src11_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src11_channel,                                                    --                .channel
			rf_sink_ready           => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                  --     (terminated)
		);

	control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                             --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                -- (terminated)
			csr_read          => '0',                                                                                 -- (terminated)
			csr_write         => '0',                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                  -- (terminated)
			almost_full_data  => open,                                                                                -- (terminated)
			almost_empty_data => open,                                                                                -- (terminated)
			in_empty          => '0',                                                                                 -- (terminated)
			out_empty         => open,                                                                                -- (terminated)
			in_error          => '0',                                                                                 -- (terminated)
			out_error         => open,                                                                                -- (terminated)
			in_channel        => '0',                                                                                 -- (terminated)
			out_channel       => open                                                                                 -- (terminated)
		);

	control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                       --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			in_data           => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_startofpacket  => '0',                                                                           -- (terminated)
			in_endofpacket    => '0',                                                                           -- (terminated)
			out_startofpacket => open,                                                                          -- (terminated)
			out_endofpacket   => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	fft_in_0_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                               --       clk_reset.reset
			m0_address              => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src12_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src12_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_002_src12_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src12_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src12_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src12_channel,                                                 --                .channel
			rf_sink_ready           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                               -- clk_reset.reset
			in_data           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                         -- clk_reset.reset
			in_data           => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                       -- (terminated)
			csr_read          => '0',                                                                        -- (terminated)
			csr_write         => '0',                                                                        -- (terminated)
			csr_readdata      => open,                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                         -- (terminated)
			almost_full_data  => open,                                                                       -- (terminated)
			almost_empty_data => open,                                                                       -- (terminated)
			in_startofpacket  => '0',                                                                        -- (terminated)
			in_endofpacket    => '0',                                                                        -- (terminated)
			out_startofpacket => open,                                                                       -- (terminated)
			out_endofpacket   => open,                                                                       -- (terminated)
			in_empty          => '0',                                                                        -- (terminated)
			out_empty         => open,                                                                       -- (terminated)
			in_error          => '0',                                                                        -- (terminated)
			out_error         => open,                                                                       -- (terminated)
			in_channel        => '0',                                                                        -- (terminated)
			out_channel       => open                                                                        -- (terminated)
		);

	fft_in_1_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                               --       clk_reset.reset
			m0_address              => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src13_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src13_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_002_src13_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src13_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src13_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src13_channel,                                                 --                .channel
			rf_sink_ready           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                               -- clk_reset.reset
			in_data           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                         -- clk_reset.reset
			in_data           => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                       -- (terminated)
			csr_read          => '0',                                                                        -- (terminated)
			csr_write         => '0',                                                                        -- (terminated)
			csr_readdata      => open,                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                         -- (terminated)
			almost_full_data  => open,                                                                       -- (terminated)
			almost_empty_data => open,                                                                       -- (terminated)
			in_startofpacket  => '0',                                                                        -- (terminated)
			in_endofpacket    => '0',                                                                        -- (terminated)
			out_startofpacket => open,                                                                       -- (terminated)
			out_endofpacket   => open,                                                                       -- (terminated)
			in_empty          => '0',                                                                        -- (terminated)
			out_empty         => open,                                                                       -- (terminated)
			in_error          => '0',                                                                        -- (terminated)
			out_error         => open,                                                                       -- (terminated)
			in_channel        => '0',                                                                        -- (terminated)
			out_channel       => open                                                                        -- (terminated)
		);

	fft_in_2_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                               --       clk_reset.reset
			m0_address              => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src14_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src14_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_002_src14_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src14_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src14_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src14_channel,                                                 --                .channel
			rf_sink_ready           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                               -- clk_reset.reset
			in_data           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                         -- clk_reset.reset
			in_data           => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                       -- (terminated)
			csr_read          => '0',                                                                        -- (terminated)
			csr_write         => '0',                                                                        -- (terminated)
			csr_readdata      => open,                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                         -- (terminated)
			almost_full_data  => open,                                                                       -- (terminated)
			almost_empty_data => open,                                                                       -- (terminated)
			in_startofpacket  => '0',                                                                        -- (terminated)
			in_endofpacket    => '0',                                                                        -- (terminated)
			out_startofpacket => open,                                                                       -- (terminated)
			out_endofpacket   => open,                                                                       -- (terminated)
			in_empty          => '0',                                                                        -- (terminated)
			out_empty         => open,                                                                       -- (terminated)
			in_error          => '0',                                                                        -- (terminated)
			out_error         => open,                                                                       -- (terminated)
			in_channel        => '0',                                                                        -- (terminated)
			out_channel       => open                                                                        -- (terminated)
		);

	fft_in_3_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                               --       clk_reset.reset
			m0_address              => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src15_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src15_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_002_src15_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src15_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src15_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src15_channel,                                                 --                .channel
			rf_sink_ready           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                               -- clk_reset.reset
			in_data           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                         -- clk_reset.reset
			in_data           => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                       -- (terminated)
			csr_read          => '0',                                                                        -- (terminated)
			csr_write         => '0',                                                                        -- (terminated)
			csr_readdata      => open,                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                         -- (terminated)
			almost_full_data  => open,                                                                       -- (terminated)
			almost_empty_data => open,                                                                       -- (terminated)
			in_startofpacket  => '0',                                                                        -- (terminated)
			in_endofpacket    => '0',                                                                        -- (terminated)
			out_startofpacket => open,                                                                       -- (terminated)
			out_endofpacket   => open,                                                                       -- (terminated)
			in_empty          => '0',                                                                        -- (terminated)
			out_empty         => open,                                                                       -- (terminated)
			in_error          => '0',                                                                        -- (terminated)
			out_error         => open,                                                                       -- (terminated)
			in_channel        => '0',                                                                        -- (terminated)
			out_channel       => open                                                                        -- (terminated)
		);

	rotary_in_s1_translator_avalon_universal_slave_0_agent : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                           --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_002_src16_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_002_src16_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_002_src16_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_002_src16_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_002_src16_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_002_src16_channel,                                                  --                .channel
			rf_sink_ready           => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                           --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                -- clk_reset.reset
			in_data           => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios2vga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			in_data           => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_startofpacket  => '0',                                                                         -- (terminated)
			in_endofpacket    => '0',                                                                         -- (terminated)
			out_startofpacket => open,                                                                        -- (terminated)
			out_endofpacket   => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	addr_router : component nios2VGA_addr_router
		port map (
			sink_ready         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                              --       src.ready
			src_valid          => addr_router_src_valid,                                                              --          .valid
			src_data           => addr_router_src_data,                                                               --          .data
			src_channel        => addr_router_src_channel,                                                            --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                         --          .endofpacket
		);

	addr_router_001 : component nios2VGA_addr_router_001
		port map (
			sink_ready         => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                                          --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                                   -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                                            --       src.ready
			src_valid          => addr_router_001_src_valid,                                                                            --          .valid
			src_data           => addr_router_001_src_data,                                                                             --          .data
			src_channel        => addr_router_001_src_channel,                                                                          --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                                    --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                                       --          .endofpacket
		);

	addr_router_002 : component nios2VGA_addr_router_002
		port map (
			sink_ready         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_002_src_ready,                                                   --       src.ready
			src_valid          => addr_router_002_src_valid,                                                   --          .valid
			src_data           => addr_router_002_src_data,                                                    --          .data
			src_channel        => addr_router_002_src_channel,                                                 --          .channel
			src_startofpacket  => addr_router_002_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => addr_router_002_src_endofpacket                                              --          .endofpacket
		);

	id_router : component nios2VGA_id_router
		port map (
			sink_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                              --       src.ready
			src_valid          => id_router_src_valid,                                                              --          .valid
			src_data           => id_router_src_data,                                                               --          .data
			src_channel        => id_router_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                         --          .endofpacket
		);

	id_router_001 : component nios2VGA_id_router_001
		port map (
			sink_ready         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                       --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                           --       src.ready
			src_valid          => id_router_001_src_valid,                                                           --          .valid
			src_data           => id_router_001_src_data,                                                            --          .data
			src_channel        => id_router_001_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                      --          .endofpacket
		);

	id_router_002 : component nios2VGA_id_router_002
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                --       src.ready
			src_valid          => id_router_002_src_valid,                                                                --          .valid
			src_data           => id_router_002_src_data,                                                                 --          .data
			src_channel        => id_router_002_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                           --          .endofpacket
		);

	id_router_003 : component nios2VGA_id_router_002
		port map (
			sink_ready         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                     --       src.ready
			src_valid          => id_router_003_src_valid,                                                     --          .valid
			src_data           => id_router_003_src_data,                                                      --          .data
			src_channel        => id_router_003_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                --          .endofpacket
		);

	id_router_004 : component nios2VGA_id_router_002
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                        --       src.ready
			src_valid          => id_router_004_src_valid,                                                        --          .valid
			src_data           => id_router_004_src_data,                                                         --          .data
			src_channel        => id_router_004_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                   --          .endofpacket
		);

	id_router_005 : component nios2VGA_id_router_002
		port map (
			sink_ready         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                   --       src.ready
			src_valid          => id_router_005_src_valid,                                                   --          .valid
			src_data           => id_router_005_src_data,                                                    --          .data
			src_channel        => id_router_005_src_channel,                                                 --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                              --          .endofpacket
		);

	id_router_006 : component nios2VGA_id_router_002
		port map (
			sink_ready         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                                               --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                                        -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                                                   --       src.ready
			src_valid          => id_router_006_src_valid,                                                                                   --          .valid
			src_data           => id_router_006_src_data,                                                                                    --          .data
			src_channel        => id_router_006_src_channel,                                                                                 --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                                           --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                                              --          .endofpacket
		);

	id_router_007 : component nios2VGA_id_router_007
		port map (
			sink_ready         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                                              --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                                       -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                                                  --       src.ready
			src_valid          => id_router_007_src_valid,                                                                                  --          .valid
			src_data           => id_router_007_src_data,                                                                                   --          .data
			src_channel        => id_router_007_src_channel,                                                                                --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                                          --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                                             --          .endofpacket
		);

	id_router_008 : component nios2VGA_id_router_002
		port map (
			sink_ready         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                                      --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                               -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                                          --       src.ready
			src_valid          => id_router_008_src_valid,                                                                          --          .valid
			src_data           => id_router_008_src_data,                                                                           --          .data
			src_channel        => id_router_008_src_channel,                                                                        --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                                                  --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                                     --          .endofpacket
		);

	id_router_009 : component nios2VGA_id_router_002
		port map (
			sink_ready         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                     --       src.ready
			src_valid          => id_router_009_src_valid,                                                     --          .valid
			src_data           => id_router_009_src_data,                                                      --          .data
			src_channel        => id_router_009_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                --          .endofpacket
		);

	id_router_010 : component nios2VGA_id_router_002
		port map (
			sink_ready         => control_in_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => control_in_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => control_in_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => control_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => control_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                  --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                                  --       src.ready
			src_valid          => id_router_010_src_valid,                                                  --          .valid
			src_data           => id_router_010_src_data,                                                   --          .data
			src_channel        => id_router_010_src_channel,                                                --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                             --          .endofpacket
		);

	id_router_011 : component nios2VGA_id_router_002
		port map (
			sink_ready         => control_out_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => control_out_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => control_out_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => control_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => control_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                   --       src.ready
			src_valid          => id_router_011_src_valid,                                                   --          .valid
			src_data           => id_router_011_src_data,                                                    --          .data
			src_channel        => id_router_011_src_channel,                                                 --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                              --          .endofpacket
		);

	id_router_012 : component nios2VGA_id_router_002
		port map (
			sink_ready         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                     -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                                --       src.ready
			src_valid          => id_router_012_src_valid,                                                --          .valid
			src_data           => id_router_012_src_data,                                                 --          .data
			src_channel        => id_router_012_src_channel,                                              --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                           --          .endofpacket
		);

	id_router_013 : component nios2VGA_id_router_002
		port map (
			sink_ready         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                     -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                                --       src.ready
			src_valid          => id_router_013_src_valid,                                                --          .valid
			src_data           => id_router_013_src_data,                                                 --          .data
			src_channel        => id_router_013_src_channel,                                              --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                           --          .endofpacket
		);

	id_router_014 : component nios2VGA_id_router_002
		port map (
			sink_ready         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                     -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                                --       src.ready
			src_valid          => id_router_014_src_valid,                                                --          .valid
			src_data           => id_router_014_src_data,                                                 --          .data
			src_channel        => id_router_014_src_channel,                                              --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                           --          .endofpacket
		);

	id_router_015 : component nios2VGA_id_router_002
		port map (
			sink_ready         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                     -- clk_reset.reset
			src_ready          => id_router_015_src_ready,                                                --       src.ready
			src_valid          => id_router_015_src_valid,                                                --          .valid
			src_data           => id_router_015_src_data,                                                 --          .data
			src_channel        => id_router_015_src_channel,                                              --          .channel
			src_startofpacket  => id_router_015_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_015_src_endofpacket                                           --          .endofpacket
		);

	id_router_016 : component nios2VGA_id_router_002
		port map (
			sink_ready         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                 --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_016_src_ready,                                                 --       src.ready
			src_valid          => id_router_016_src_valid,                                                 --          .valid
			src_data           => id_router_016_src_data,                                                  --          .data
			src_channel        => id_router_016_src_channel,                                               --          .channel
			src_startofpacket  => id_router_016_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_016_src_endofpacket                                            --          .endofpacket
		);

	burst_adapter : component nios2vga_burst_adapter
		generic map (
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 69,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 64,
			PKT_BURST_SIZE_L          => 62,
			PKT_BURST_TYPE_H          => 66,
			PKT_BURST_TYPE_L          => 65,
			PKT_BURSTWRAP_H           => 61,
			PKT_BURSTWRAP_L           => 59,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 91,
			ST_CHANNEL_W              => 17,
			OUT_BYTE_CNT_H            => 57,
			OUT_BURSTWRAP_H           => 61,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => external_clocks_sys_clk_clk,         --       cr0.clk
			reset                 => rst_controller_002_reset_out_reset,  -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_001_src_valid,          --     sink0.valid
			sink0_data            => cmd_xbar_mux_001_src_data,           --          .data
			sink0_channel         => cmd_xbar_mux_001_src_channel,        --          .channel
			sink0_startofpacket   => cmd_xbar_mux_001_src_startofpacket,  --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_001_src_endofpacket,    --          .endofpacket
			sink0_ready           => cmd_xbar_mux_001_src_ready,          --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component nios2vga_burst_adapter_001
		generic map (
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_BEGIN_BURST           => 60,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_BURST_SIZE_H          => 55,
			PKT_BURST_SIZE_L          => 53,
			PKT_BURST_TYPE_H          => 57,
			PKT_BURST_TYPE_L          => 56,
			PKT_BURSTWRAP_H           => 52,
			PKT_BURSTWRAP_L           => 50,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 82,
			ST_CHANNEL_W              => 17,
			OUT_BYTE_CNT_H            => 47,
			OUT_BURSTWRAP_H           => 52,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 7,
			BURSTWRAP_CONST_VALUE     => 7
		)
		port map (
			clk                   => external_clocks_sys_clk_clk,             --       cr0.clk
			reset                 => rst_controller_002_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => crosser_006_out_valid,                   --     sink0.valid
			sink0_data            => crosser_006_out_data,                    --          .data
			sink0_channel         => crosser_006_out_channel,                 --          .channel
			sink0_startofpacket   => crosser_006_out_startofpacket,           --          .startofpacket
			sink0_endofpacket     => crosser_006_out_endofpacket,             --          .endofpacket
			sink0_ready           => crosser_006_out_ready,                   --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	rst_controller : component nios2vga_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,                       -- reset_in0.reset
			reset_in1  => external_clocks_sys_clk_reset_reset_ports_inv, -- reset_in1.reset
			clk        => clk_clk,                                       --       clk.clk
			reset_out  => rst_controller_reset_out_reset,                -- reset_out.reset
			reset_req  => open,                                          -- (terminated)
			reset_in2  => '0',                                           -- (terminated)
			reset_in3  => '0',                                           -- (terminated)
			reset_in4  => '0',                                           -- (terminated)
			reset_in5  => '0',                                           -- (terminated)
			reset_in6  => '0',                                           -- (terminated)
			reset_in7  => '0',                                           -- (terminated)
			reset_in8  => '0',                                           -- (terminated)
			reset_in9  => '0',                                           -- (terminated)
			reset_in10 => '0',                                           -- (terminated)
			reset_in11 => '0',                                           -- (terminated)
			reset_in12 => '0',                                           -- (terminated)
			reset_in13 => '0',                                           -- (terminated)
			reset_in14 => '0',                                           -- (terminated)
			reset_in15 => '0'                                            -- (terminated)
		);

	rst_controller_001 : component nios2vga_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => clk_clk,                            --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component nios2vga_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset,  -- reset_in1.reset
			clk        => external_clocks_sys_clk_clk,        --       clk.clk
			reset_out  => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component nios2vga_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset,  -- reset_in1.reset
			clk        => external_clocks_vga_clk_clk,        --       clk.clk
			reset_out  => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component nios2VGA_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component nios2VGA_cmd_xbar_demux_001
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_001_src_ready,             --      sink.ready
			sink_channel       => addr_router_001_src_channel,           --          .channel
			sink_data          => addr_router_001_src_data,              --          .data
			sink_startofpacket => addr_router_001_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_001_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_001_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_002 : component nios2VGA_cmd_xbar_demux_002
		port map (
			clk                 => clk_clk,                                --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			sink_ready          => addr_router_002_src_ready,              --      sink.ready
			sink_channel        => addr_router_002_src_channel,            --          .channel
			sink_data           => addr_router_002_src_data,               --          .data
			sink_startofpacket  => addr_router_002_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_002_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_002_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_002_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_002_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_002_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_002_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_002_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_002_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_002_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_002_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_002_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_002_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_002_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_002_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_002_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_002_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_002_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_002_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_002_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_002_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_002_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_002_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_002_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_002_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_002_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_002_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_002_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_002_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_002_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_002_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_002_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_002_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_002_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_002_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_002_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_002_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_002_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_002_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_002_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_002_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_002_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_002_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_002_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_002_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_002_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_002_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_002_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_002_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_002_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_002_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_002_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_002_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_002_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_002_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_002_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_002_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_002_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_002_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_002_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_002_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_002_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_002_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_002_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_002_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_002_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_002_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_002_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_002_src10_endofpacket,   --          .endofpacket
			src11_ready         => cmd_xbar_demux_002_src11_ready,         --     src11.ready
			src11_valid         => cmd_xbar_demux_002_src11_valid,         --          .valid
			src11_data          => cmd_xbar_demux_002_src11_data,          --          .data
			src11_channel       => cmd_xbar_demux_002_src11_channel,       --          .channel
			src11_startofpacket => cmd_xbar_demux_002_src11_startofpacket, --          .startofpacket
			src11_endofpacket   => cmd_xbar_demux_002_src11_endofpacket,   --          .endofpacket
			src12_ready         => cmd_xbar_demux_002_src12_ready,         --     src12.ready
			src12_valid         => cmd_xbar_demux_002_src12_valid,         --          .valid
			src12_data          => cmd_xbar_demux_002_src12_data,          --          .data
			src12_channel       => cmd_xbar_demux_002_src12_channel,       --          .channel
			src12_startofpacket => cmd_xbar_demux_002_src12_startofpacket, --          .startofpacket
			src12_endofpacket   => cmd_xbar_demux_002_src12_endofpacket,   --          .endofpacket
			src13_ready         => cmd_xbar_demux_002_src13_ready,         --     src13.ready
			src13_valid         => cmd_xbar_demux_002_src13_valid,         --          .valid
			src13_data          => cmd_xbar_demux_002_src13_data,          --          .data
			src13_channel       => cmd_xbar_demux_002_src13_channel,       --          .channel
			src13_startofpacket => cmd_xbar_demux_002_src13_startofpacket, --          .startofpacket
			src13_endofpacket   => cmd_xbar_demux_002_src13_endofpacket,   --          .endofpacket
			src14_ready         => cmd_xbar_demux_002_src14_ready,         --     src14.ready
			src14_valid         => cmd_xbar_demux_002_src14_valid,         --          .valid
			src14_data          => cmd_xbar_demux_002_src14_data,          --          .data
			src14_channel       => cmd_xbar_demux_002_src14_channel,       --          .channel
			src14_startofpacket => cmd_xbar_demux_002_src14_startofpacket, --          .startofpacket
			src14_endofpacket   => cmd_xbar_demux_002_src14_endofpacket,   --          .endofpacket
			src15_ready         => cmd_xbar_demux_002_src15_ready,         --     src15.ready
			src15_valid         => cmd_xbar_demux_002_src15_valid,         --          .valid
			src15_data          => cmd_xbar_demux_002_src15_data,          --          .data
			src15_channel       => cmd_xbar_demux_002_src15_channel,       --          .channel
			src15_startofpacket => cmd_xbar_demux_002_src15_startofpacket, --          .startofpacket
			src15_endofpacket   => cmd_xbar_demux_002_src15_endofpacket,   --          .endofpacket
			src16_ready         => cmd_xbar_demux_002_src16_ready,         --     src16.ready
			src16_valid         => cmd_xbar_demux_002_src16_valid,         --          .valid
			src16_data          => cmd_xbar_demux_002_src16_data,          --          .data
			src16_channel       => cmd_xbar_demux_002_src16_channel,       --          .channel
			src16_startofpacket => cmd_xbar_demux_002_src16_startofpacket, --          .startofpacket
			src16_endofpacket   => cmd_xbar_demux_002_src16_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component nios2VGA_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_002_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_002_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component nios2VGA_cmd_xbar_mux_001
		port map (
			clk                 => external_clocks_sys_clk_clk,           --       clk.clk
			reset               => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => crosser_004_out_ready,                 --     sink0.ready
			sink0_valid         => crosser_004_out_valid,                 --          .valid
			sink0_channel       => crosser_004_out_channel,               --          .channel
			sink0_data          => crosser_004_out_data,                  --          .data
			sink0_startofpacket => crosser_004_out_startofpacket,         --          .startofpacket
			sink0_endofpacket   => crosser_004_out_endofpacket,           --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => crosser_005_out_ready,                 --     sink2.ready
			sink2_valid         => crosser_005_out_valid,                 --          .valid
			sink2_channel       => crosser_005_out_channel,               --          .channel
			sink2_data          => crosser_005_out_data,                  --          .data
			sink2_startofpacket => crosser_005_out_startofpacket,         --          .startofpacket
			sink2_endofpacket   => crosser_005_out_endofpacket            --          .endofpacket
		);

	rsp_xbar_demux : component nios2VGA_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component nios2VGA_rsp_xbar_demux_001
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			src2_ready         => rsp_xbar_demux_001_src2_ready,         --      src2.ready
			src2_valid         => rsp_xbar_demux_001_src2_valid,         --          .valid
			src2_data          => rsp_xbar_demux_001_src2_data,          --          .data
			src2_channel       => rsp_xbar_demux_001_src2_channel,       --          .channel
			src2_startofpacket => rsp_xbar_demux_001_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => rsp_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component nios2VGA_rsp_xbar_demux_007
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_014_src_ready,               --      sink.ready
			sink_channel       => id_router_014_src_channel,             --          .channel
			sink_data          => id_router_014_src_data,                --          .data
			sink_startofpacket => id_router_014_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_014_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_014_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_015 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_015_src_ready,               --      sink.ready
			sink_channel       => id_router_015_src_channel,             --          .channel
			sink_data          => id_router_015_src_data,                --          .data
			sink_startofpacket => id_router_015_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_015_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_015_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_015_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_015_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_015_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_016 : component nios2VGA_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_016_src_ready,               --      sink.ready
			sink_channel       => id_router_016_src_channel,             --          .channel
			sink_data          => id_router_016_src_data,                --          .data
			sink_startofpacket => id_router_016_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_016_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_016_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_016_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_016_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_016_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component nios2VGA_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,    -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_src_data,             --          .data
			src_channel         => rsp_xbar_mux_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,         --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,          --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			sink1_ready         => crosser_007_out_ready,             --     sink1.ready
			sink1_valid         => crosser_007_out_valid,             --          .valid
			sink1_channel       => crosser_007_out_channel,           --          .channel
			sink1_data          => crosser_007_out_data,              --          .data
			sink1_startofpacket => crosser_007_out_startofpacket,     --          .startofpacket
			sink1_endofpacket   => crosser_007_out_endofpacket        --          .endofpacket
		);

	rsp_xbar_mux_002 : component nios2VGA_rsp_xbar_mux_002
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_002_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_002_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_002_src_data,             --          .data
			src_channel          => rsp_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => crosser_008_out_ready,                 --     sink1.ready
			sink1_valid          => crosser_008_out_valid,                 --          .valid
			sink1_channel        => crosser_008_out_channel,               --          .channel
			sink1_data           => crosser_008_out_data,                  --          .data
			sink1_startofpacket  => crosser_008_out_startofpacket,         --          .startofpacket
			sink1_endofpacket    => crosser_008_out_endofpacket,           --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => crosser_002_out_ready,                 --     sink6.ready
			sink6_valid          => crosser_002_out_valid,                 --          .valid
			sink6_channel        => crosser_002_out_channel,               --          .channel
			sink6_data           => crosser_002_out_data,                  --          .data
			sink6_startofpacket  => crosser_002_out_startofpacket,         --          .startofpacket
			sink6_endofpacket    => crosser_002_out_endofpacket,           --          .endofpacket
			sink7_ready          => crosser_009_out_ready,                 --     sink7.ready
			sink7_valid          => crosser_009_out_valid,                 --          .valid
			sink7_channel        => crosser_009_out_channel,               --          .channel
			sink7_data           => crosser_009_out_data,                  --          .data
			sink7_startofpacket  => crosser_009_out_startofpacket,         --          .startofpacket
			sink7_endofpacket    => crosser_009_out_endofpacket,           --          .endofpacket
			sink8_ready          => crosser_003_out_ready,                 --     sink8.ready
			sink8_valid          => crosser_003_out_valid,                 --          .valid
			sink8_channel        => crosser_003_out_channel,               --          .channel
			sink8_data           => crosser_003_out_data,                  --          .data
			sink8_startofpacket  => crosser_003_out_startofpacket,         --          .startofpacket
			sink8_endofpacket    => crosser_003_out_endofpacket,           --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink14_ready         => rsp_xbar_demux_014_src0_ready,         --    sink14.ready
			sink14_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink14_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink14_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink14_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink14_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			sink15_ready         => rsp_xbar_demux_015_src0_ready,         --    sink15.ready
			sink15_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			sink15_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			sink15_data          => rsp_xbar_demux_015_src0_data,          --          .data
			sink15_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			sink15_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			sink16_ready         => rsp_xbar_demux_016_src0_ready,         --    sink16.ready
			sink16_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			sink16_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			sink16_data          => rsp_xbar_demux_016_src0_data,          --          .data
			sink16_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			sink16_endofpacket   => rsp_xbar_demux_016_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component nios2vga_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 79,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 82,
			IN_PKT_BURST_SIZE_L           => 80,
			IN_PKT_RESPONSE_STATUS_H      => 108,
			IN_PKT_RESPONSE_STATUS_L      => 107,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 84,
			IN_PKT_BURST_TYPE_L           => 83,
			IN_ST_DATA_W                  => 109,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 58,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 64,
			OUT_PKT_BURST_SIZE_L          => 62,
			OUT_PKT_RESPONSE_STATUS_H     => 90,
			OUT_PKT_RESPONSE_STATUS_L     => 89,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 66,
			OUT_PKT_BURST_TYPE_L          => 65,
			OUT_ST_DATA_W                 => 91,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                           --       clk.clk
			reset                => rst_controller_reset_out_reset,    -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src1_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_src1_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src1_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_src1_ready,         --          .ready
			in_data              => cmd_xbar_demux_src1_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_src_data,            --          .data
			out_channel          => width_adapter_src_channel,         --          .channel
			out_valid            => width_adapter_src_valid,           --          .valid
			out_ready            => width_adapter_src_ready,           --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                              -- (terminated)
		);

	width_adapter_001 : component nios2vga_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 79,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 82,
			IN_PKT_BURST_SIZE_L           => 80,
			IN_PKT_RESPONSE_STATUS_H      => 108,
			IN_PKT_RESPONSE_STATUS_L      => 107,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 84,
			IN_PKT_BURST_TYPE_L           => 83,
			IN_ST_DATA_W                  => 109,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 58,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 64,
			OUT_PKT_BURST_SIZE_L          => 62,
			OUT_PKT_RESPONSE_STATUS_H     => 90,
			OUT_PKT_RESPONSE_STATUS_L     => 89,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 66,
			OUT_PKT_BURST_TYPE_L          => 65,
			OUT_ST_DATA_W                 => 91,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_002_src1_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_002_src1_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_002_src1_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_002_src1_ready,         --          .ready
			in_data              => cmd_xbar_demux_002_src1_data,          --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_001_src_data,            --          .data
			out_channel          => width_adapter_001_src_channel,         --          .channel
			out_valid            => width_adapter_001_src_valid,           --          .valid
			out_ready            => width_adapter_001_src_ready,           --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_002 : component nios2vga_width_adapter_002
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 79,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 82,
			IN_PKT_BURST_SIZE_L           => 80,
			IN_PKT_RESPONSE_STATUS_H      => 108,
			IN_PKT_RESPONSE_STATUS_L      => 107,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 84,
			IN_PKT_BURST_TYPE_L           => 83,
			IN_ST_DATA_W                  => 109,
			OUT_PKT_ADDR_H                => 40,
			OUT_PKT_ADDR_L                => 9,
			OUT_PKT_DATA_H                => 7,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 8,
			OUT_PKT_BYTEEN_L              => 8,
			OUT_PKT_BYTE_CNT_H            => 49,
			OUT_PKT_BYTE_CNT_L            => 47,
			OUT_PKT_TRANS_COMPRESSED_READ => 41,
			OUT_PKT_BURST_SIZE_H          => 55,
			OUT_PKT_BURST_SIZE_L          => 53,
			OUT_PKT_RESPONSE_STATUS_H     => 81,
			OUT_PKT_RESPONSE_STATUS_L     => 80,
			OUT_PKT_TRANS_EXCLUSIVE       => 46,
			OUT_PKT_BURST_TYPE_H          => 57,
			OUT_PKT_BURST_TYPE_L          => 56,
			OUT_ST_DATA_W                 => 82,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_002_src7_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_002_src7_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_002_src7_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_002_src7_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_002_src7_ready,         --          .ready
			in_data              => cmd_xbar_demux_002_src7_data,          --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_002_src_data,            --          .data
			out_channel          => width_adapter_002_src_channel,         --          .channel
			out_valid            => width_adapter_002_src_valid,           --          .valid
			out_ready            => width_adapter_002_src_ready,           --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_003 : component nios2vga_width_adapter_003
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 58,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 61,
			IN_PKT_BURSTWRAP_L            => 59,
			IN_PKT_BURST_SIZE_H           => 64,
			IN_PKT_BURST_SIZE_L           => 62,
			IN_PKT_RESPONSE_STATUS_H      => 90,
			IN_PKT_RESPONSE_STATUS_L      => 89,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 66,
			IN_PKT_BURST_TYPE_L           => 65,
			IN_ST_DATA_W                  => 91,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 82,
			OUT_PKT_BURST_SIZE_L          => 80,
			OUT_PKT_RESPONSE_STATUS_H     => 108,
			OUT_PKT_RESPONSE_STATUS_L     => 107,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 84,
			OUT_PKT_BURST_TYPE_L          => 83,
			OUT_ST_DATA_W                 => 109,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => external_clocks_sys_clk_clk,           --       clk.clk
			reset                => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			in_valid             => rsp_xbar_demux_001_src0_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_001_src0_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_001_src0_ready,         --          .ready
			in_data              => rsp_xbar_demux_001_src0_data,          --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_003_src_data,            --          .data
			out_channel          => width_adapter_003_src_channel,         --          .channel
			out_valid            => width_adapter_003_src_valid,           --          .valid
			out_ready            => width_adapter_003_src_ready,           --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_004 : component nios2vga_width_adapter_003
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 58,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 61,
			IN_PKT_BURSTWRAP_L            => 59,
			IN_PKT_BURST_SIZE_H           => 64,
			IN_PKT_BURST_SIZE_L           => 62,
			IN_PKT_RESPONSE_STATUS_H      => 90,
			IN_PKT_RESPONSE_STATUS_L      => 89,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 66,
			IN_PKT_BURST_TYPE_L           => 65,
			IN_ST_DATA_W                  => 91,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 82,
			OUT_PKT_BURST_SIZE_L          => 80,
			OUT_PKT_RESPONSE_STATUS_H     => 108,
			OUT_PKT_RESPONSE_STATUS_L     => 107,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 84,
			OUT_PKT_BURST_TYPE_L          => 83,
			OUT_ST_DATA_W                 => 109,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => external_clocks_sys_clk_clk,           --       clk.clk
			reset                => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			in_valid             => rsp_xbar_demux_001_src2_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_001_src2_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_001_src2_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_001_src2_ready,         --          .ready
			in_data              => rsp_xbar_demux_001_src2_data,          --          .data
			out_endofpacket      => width_adapter_004_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_004_src_data,            --          .data
			out_channel          => width_adapter_004_src_channel,         --          .channel
			out_valid            => width_adapter_004_src_valid,           --          .valid
			out_ready            => width_adapter_004_src_ready,           --          .ready
			out_startofpacket    => width_adapter_004_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_005 : component nios2vga_width_adapter_005
		generic map (
			IN_PKT_ADDR_H                 => 40,
			IN_PKT_ADDR_L                 => 9,
			IN_PKT_DATA_H                 => 7,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 8,
			IN_PKT_BYTEEN_L               => 8,
			IN_PKT_BYTE_CNT_H             => 49,
			IN_PKT_BYTE_CNT_L             => 47,
			IN_PKT_TRANS_COMPRESSED_READ  => 41,
			IN_PKT_BURSTWRAP_H            => 52,
			IN_PKT_BURSTWRAP_L            => 50,
			IN_PKT_BURST_SIZE_H           => 55,
			IN_PKT_BURST_SIZE_L           => 53,
			IN_PKT_RESPONSE_STATUS_H      => 81,
			IN_PKT_RESPONSE_STATUS_L      => 80,
			IN_PKT_TRANS_EXCLUSIVE        => 46,
			IN_PKT_BURST_TYPE_H           => 57,
			IN_PKT_BURST_TYPE_L           => 56,
			IN_ST_DATA_W                  => 82,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 82,
			OUT_PKT_BURST_SIZE_L          => 80,
			OUT_PKT_RESPONSE_STATUS_H     => 108,
			OUT_PKT_RESPONSE_STATUS_L     => 107,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 84,
			OUT_PKT_BURST_TYPE_L          => 83,
			OUT_ST_DATA_W                 => 109,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => external_clocks_sys_clk_clk,           --       clk.clk
			reset                => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			in_valid             => rsp_xbar_demux_007_src0_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_007_src0_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_007_src0_ready,         --          .ready
			in_data              => rsp_xbar_demux_007_src0_data,          --          .data
			out_endofpacket      => width_adapter_005_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_005_src_data,            --          .data
			out_channel          => width_adapter_005_src_channel,         --          .channel
			out_valid            => width_adapter_005_src_valid,           --          .valid
			out_ready            => width_adapter_005_src_ready,           --          .ready
			out_startofpacket    => width_adapter_005_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	crosser : component nios2vga_crosser
		generic map (
			DATA_WIDTH          => 109,
			BITS_PER_SYMBOL     => 109,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => external_clocks_sys_clk_clk,           --       out_clk.clk
			out_reset         => rst_controller_002_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src6_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src6_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src6_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src6_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src6_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src6_data,          --              .data
			out_ready         => crosser_out_ready,                     --           out.ready
			out_valid         => crosser_out_valid,                     --              .valid
			out_startofpacket => crosser_out_startofpacket,             --              .startofpacket
			out_endofpacket   => crosser_out_endofpacket,               --              .endofpacket
			out_channel       => crosser_out_channel,                   --              .channel
			out_data          => crosser_out_data,                      --              .data
			in_empty          => '0',                                   --   (terminated)
			in_error          => '0',                                   --   (terminated)
			out_empty         => open,                                  --   (terminated)
			out_error         => open                                   --   (terminated)
		);

	crosser_001 : component nios2vga_crosser
		generic map (
			DATA_WIDTH          => 109,
			BITS_PER_SYMBOL     => 109,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => clk_clk,                               --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => external_clocks_sys_clk_clk,           --       out_clk.clk
			out_reset         => rst_controller_002_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_002_src8_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_002_src8_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_002_src8_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_002_src8_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_002_src8_channel,       --              .channel
			in_data           => cmd_xbar_demux_002_src8_data,          --              .data
			out_ready         => crosser_001_out_ready,                 --           out.ready
			out_valid         => crosser_001_out_valid,                 --              .valid
			out_startofpacket => crosser_001_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_001_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_001_out_channel,               --              .channel
			out_data          => crosser_001_out_data,                  --              .data
			in_empty          => '0',                                   --   (terminated)
			in_error          => '0',                                   --   (terminated)
			out_empty         => open,                                  --   (terminated)
			out_error         => open                                   --   (terminated)
		);

	crosser_002 : component nios2vga_crosser
		generic map (
			DATA_WIDTH          => 109,
			BITS_PER_SYMBOL     => 109,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => external_clocks_sys_clk_clk,           --        in_clk.clk
			in_reset          => rst_controller_002_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_006_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_006_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_006_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_006_src0_data,          --              .data
			out_ready         => crosser_002_out_ready,                 --           out.ready
			out_valid         => crosser_002_out_valid,                 --              .valid
			out_startofpacket => crosser_002_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_002_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_002_out_channel,               --              .channel
			out_data          => crosser_002_out_data,                  --              .data
			in_empty          => '0',                                   --   (terminated)
			in_error          => '0',                                   --   (terminated)
			out_empty         => open,                                  --   (terminated)
			out_error         => open                                   --   (terminated)
		);

	crosser_003 : component nios2vga_crosser
		generic map (
			DATA_WIDTH          => 109,
			BITS_PER_SYMBOL     => 109,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => external_clocks_sys_clk_clk,           --        in_clk.clk
			in_reset          => rst_controller_002_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => clk_clk,                               --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_008_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_008_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_008_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_008_src0_data,          --              .data
			out_ready         => crosser_003_out_ready,                 --           out.ready
			out_valid         => crosser_003_out_valid,                 --              .valid
			out_startofpacket => crosser_003_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_003_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_003_out_channel,               --              .channel
			out_data          => crosser_003_out_data,                  --              .data
			in_empty          => '0',                                   --   (terminated)
			in_error          => '0',                                   --   (terminated)
			out_empty         => open,                                  --   (terminated)
			out_error         => open                                   --   (terminated)
		);

	crosser_004 : component nios2vga_crosser_004
		generic map (
			DATA_WIDTH          => 91,
			BITS_PER_SYMBOL     => 91,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => clk_clk,                            --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,     --  in_clk_reset.reset
			out_clk           => external_clocks_sys_clk_clk,        --       out_clk.clk
			out_reset         => rst_controller_002_reset_out_reset, -- out_clk_reset.reset
			in_ready          => width_adapter_src_ready,            --            in.ready
			in_valid          => width_adapter_src_valid,            --              .valid
			in_startofpacket  => width_adapter_src_startofpacket,    --              .startofpacket
			in_endofpacket    => width_adapter_src_endofpacket,      --              .endofpacket
			in_channel        => width_adapter_src_channel,          --              .channel
			in_data           => width_adapter_src_data,             --              .data
			out_ready         => crosser_004_out_ready,              --           out.ready
			out_valid         => crosser_004_out_valid,              --              .valid
			out_startofpacket => crosser_004_out_startofpacket,      --              .startofpacket
			out_endofpacket   => crosser_004_out_endofpacket,        --              .endofpacket
			out_channel       => crosser_004_out_channel,            --              .channel
			out_data          => crosser_004_out_data,               --              .data
			in_empty          => '0',                                --   (terminated)
			in_error          => '0',                                --   (terminated)
			out_empty         => open,                               --   (terminated)
			out_error         => open                                --   (terminated)
		);

	crosser_005 : component nios2vga_crosser_004
		generic map (
			DATA_WIDTH          => 91,
			BITS_PER_SYMBOL     => 91,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => clk_clk,                             --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,      --  in_clk_reset.reset
			out_clk           => external_clocks_sys_clk_clk,         --       out_clk.clk
			out_reset         => rst_controller_002_reset_out_reset,  -- out_clk_reset.reset
			in_ready          => width_adapter_001_src_ready,         --            in.ready
			in_valid          => width_adapter_001_src_valid,         --              .valid
			in_startofpacket  => width_adapter_001_src_startofpacket, --              .startofpacket
			in_endofpacket    => width_adapter_001_src_endofpacket,   --              .endofpacket
			in_channel        => width_adapter_001_src_channel,       --              .channel
			in_data           => width_adapter_001_src_data,          --              .data
			out_ready         => crosser_005_out_ready,               --           out.ready
			out_valid         => crosser_005_out_valid,               --              .valid
			out_startofpacket => crosser_005_out_startofpacket,       --              .startofpacket
			out_endofpacket   => crosser_005_out_endofpacket,         --              .endofpacket
			out_channel       => crosser_005_out_channel,             --              .channel
			out_data          => crosser_005_out_data,                --              .data
			in_empty          => '0',                                 --   (terminated)
			in_error          => '0',                                 --   (terminated)
			out_empty         => open,                                --   (terminated)
			out_error         => open                                 --   (terminated)
		);

	crosser_006 : component nios2vga_crosser_006
		generic map (
			DATA_WIDTH          => 82,
			BITS_PER_SYMBOL     => 82,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => clk_clk,                             --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,      --  in_clk_reset.reset
			out_clk           => external_clocks_sys_clk_clk,         --       out_clk.clk
			out_reset         => rst_controller_002_reset_out_reset,  -- out_clk_reset.reset
			in_ready          => width_adapter_002_src_ready,         --            in.ready
			in_valid          => width_adapter_002_src_valid,         --              .valid
			in_startofpacket  => width_adapter_002_src_startofpacket, --              .startofpacket
			in_endofpacket    => width_adapter_002_src_endofpacket,   --              .endofpacket
			in_channel        => width_adapter_002_src_channel,       --              .channel
			in_data           => width_adapter_002_src_data,          --              .data
			out_ready         => crosser_006_out_ready,               --           out.ready
			out_valid         => crosser_006_out_valid,               --              .valid
			out_startofpacket => crosser_006_out_startofpacket,       --              .startofpacket
			out_endofpacket   => crosser_006_out_endofpacket,         --              .endofpacket
			out_channel       => crosser_006_out_channel,             --              .channel
			out_data          => crosser_006_out_data,                --              .data
			in_empty          => '0',                                 --   (terminated)
			in_error          => '0',                                 --   (terminated)
			out_empty         => open,                                --   (terminated)
			out_error         => open                                 --   (terminated)
		);

	crosser_007 : component nios2vga_crosser
		generic map (
			DATA_WIDTH          => 109,
			BITS_PER_SYMBOL     => 109,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => external_clocks_sys_clk_clk,         --        in_clk.clk
			in_reset          => rst_controller_002_reset_out_reset,  --  in_clk_reset.reset
			out_clk           => clk_clk,                             --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,      -- out_clk_reset.reset
			in_ready          => width_adapter_003_src_ready,         --            in.ready
			in_valid          => width_adapter_003_src_valid,         --              .valid
			in_startofpacket  => width_adapter_003_src_startofpacket, --              .startofpacket
			in_endofpacket    => width_adapter_003_src_endofpacket,   --              .endofpacket
			in_channel        => width_adapter_003_src_channel,       --              .channel
			in_data           => width_adapter_003_src_data,          --              .data
			out_ready         => crosser_007_out_ready,               --           out.ready
			out_valid         => crosser_007_out_valid,               --              .valid
			out_startofpacket => crosser_007_out_startofpacket,       --              .startofpacket
			out_endofpacket   => crosser_007_out_endofpacket,         --              .endofpacket
			out_channel       => crosser_007_out_channel,             --              .channel
			out_data          => crosser_007_out_data,                --              .data
			in_empty          => '0',                                 --   (terminated)
			in_error          => '0',                                 --   (terminated)
			out_empty         => open,                                --   (terminated)
			out_error         => open                                 --   (terminated)
		);

	crosser_008 : component nios2vga_crosser
		generic map (
			DATA_WIDTH          => 109,
			BITS_PER_SYMBOL     => 109,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => external_clocks_sys_clk_clk,         --        in_clk.clk
			in_reset          => rst_controller_002_reset_out_reset,  --  in_clk_reset.reset
			out_clk           => clk_clk,                             --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,      -- out_clk_reset.reset
			in_ready          => width_adapter_004_src_ready,         --            in.ready
			in_valid          => width_adapter_004_src_valid,         --              .valid
			in_startofpacket  => width_adapter_004_src_startofpacket, --              .startofpacket
			in_endofpacket    => width_adapter_004_src_endofpacket,   --              .endofpacket
			in_channel        => width_adapter_004_src_channel,       --              .channel
			in_data           => width_adapter_004_src_data,          --              .data
			out_ready         => crosser_008_out_ready,               --           out.ready
			out_valid         => crosser_008_out_valid,               --              .valid
			out_startofpacket => crosser_008_out_startofpacket,       --              .startofpacket
			out_endofpacket   => crosser_008_out_endofpacket,         --              .endofpacket
			out_channel       => crosser_008_out_channel,             --              .channel
			out_data          => crosser_008_out_data,                --              .data
			in_empty          => '0',                                 --   (terminated)
			in_error          => '0',                                 --   (terminated)
			out_empty         => open,                                --   (terminated)
			out_error         => open                                 --   (terminated)
		);

	crosser_009 : component nios2vga_crosser
		generic map (
			DATA_WIDTH          => 109,
			BITS_PER_SYMBOL     => 109,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 17,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => external_clocks_sys_clk_clk,         --        in_clk.clk
			in_reset          => rst_controller_002_reset_out_reset,  --  in_clk_reset.reset
			out_clk           => clk_clk,                             --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,      -- out_clk_reset.reset
			in_ready          => width_adapter_005_src_ready,         --            in.ready
			in_valid          => width_adapter_005_src_valid,         --              .valid
			in_startofpacket  => width_adapter_005_src_startofpacket, --              .startofpacket
			in_endofpacket    => width_adapter_005_src_endofpacket,   --              .endofpacket
			in_channel        => width_adapter_005_src_channel,       --              .channel
			in_data           => width_adapter_005_src_data,          --              .data
			out_ready         => crosser_009_out_ready,               --           out.ready
			out_valid         => crosser_009_out_valid,               --              .valid
			out_startofpacket => crosser_009_out_startofpacket,       --              .startofpacket
			out_endofpacket   => crosser_009_out_endofpacket,         --              .endofpacket
			out_channel       => crosser_009_out_channel,             --              .channel
			out_data          => crosser_009_out_data,                --              .data
			in_empty          => '0',                                 --   (terminated)
			in_error          => '0',                                 --   (terminated)
			out_empty         => open,                                --   (terminated)
			out_error         => open                                 --   (terminated)
		);

	irq_mapper : component nios2VGA_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	sys_clk_timer_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sys_clk_timer_s1_translator_avalon_anti_slave_0_write;

	red_led_pio_s1_translator_avalon_anti_slave_0_write_ports_inv <= not red_led_pio_s1_translator_avalon_anti_slave_0_write;

	green_led_pio_s1_translator_avalon_anti_slave_0_write_ports_inv <= not green_led_pio_s1_translator_avalon_anti_slave_0_write;

	control_out_s1_translator_avalon_anti_slave_0_write_ports_inv <= not control_out_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	external_clocks_sys_clk_reset_reset_ports_inv <= not external_clocks_sys_clk_reset_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	vga_clock_out_clk_clk <= external_clocks_vga_clk_clk;

end architecture rtl; -- of nios2VGA
