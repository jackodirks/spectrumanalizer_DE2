library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

ENTITY adc_sample_grabber IS
	PORT (
	ADC:    		inout std_logic_vector(11 downto 0);
	samples:   out std_logic_vector(20479 DOWNTO 0);
	clk, grab : IN std_logic;
	done : OUT STD_logic;
	sample_count : IN STD_logic_VECTOR (11 DOWNTO 0)
);
END adc_sample_grabber;

ARCHITECTURE adc_grabber OF adc_sample_grabber IS
BEGIN
	PROCESS(clk,grab,adc)
	variable temp: std_logic_vector(20479 downto 0) := (OTHERS => '0');
	BEGIN
	IF RISING_EDGE(clk) THEN
		IF (GRAB = '1') THEN
			case to_integer(unsigned(sample_count)) is
			WHEN 0 => temp(9 DOWNTO 0) := ADC(11 DOWNTO 2);
			WHEN 1 => temp(19 DOWNTO 10) := ADC(11 DOWNTO 2);
			WHEN 2 => temp(29 DOWNTO 20) := ADC(11 DOWNTO 2);
			WHEN 3 => temp(39 DOWNTO 30) := ADC(11 DOWNTO 2);
			WHEN 4 => temp(49 DOWNTO 40) := ADC(11 DOWNTO 2);
			WHEN 5 => temp(59 DOWNTO 50) := ADC(11 DOWNTO 2);
			WHEN 6 => temp(69 DOWNTO 60) := ADC(11 DOWNTO 2);
			WHEN 7 => temp(79 DOWNTO 70) := ADC(11 DOWNTO 2);
			WHEN 8 => temp(89 DOWNTO 80) := ADC(11 DOWNTO 2);
			WHEN 9 => temp(99 DOWNTO 90) := ADC(11 DOWNTO 2);
			WHEN 10 => temp(109 DOWNTO 100) := ADC(11 DOWNTO 2);
			WHEN 11 => temp(119 DOWNTO 110) := ADC(11 DOWNTO 2);
			WHEN 12 => temp(129 DOWNTO 120) := ADC(11 DOWNTO 2);
			WHEN 13 => temp(139 DOWNTO 130) := ADC(11 DOWNTO 2);
			WHEN 14 => temp(149 DOWNTO 140) := ADC(11 DOWNTO 2);
			WHEN 15 => temp(159 DOWNTO 150) := ADC(11 DOWNTO 2);
			WHEN 16 => temp(169 DOWNTO 160) := ADC(11 DOWNTO 2);
			WHEN 17 => temp(179 DOWNTO 170) := ADC(11 DOWNTO 2);
			WHEN 18 => temp(189 DOWNTO 180) := ADC(11 DOWNTO 2);
			WHEN 19 => temp(199 DOWNTO 190) := ADC(11 DOWNTO 2);
			WHEN 20 => temp(209 DOWNTO 200) := ADC(11 DOWNTO 2);
			WHEN 21 => temp(219 DOWNTO 210) := ADC(11 DOWNTO 2);
			WHEN 22 => temp(229 DOWNTO 220) := ADC(11 DOWNTO 2);
			WHEN 23 => temp(239 DOWNTO 230) := ADC(11 DOWNTO 2);
			WHEN 24 => temp(249 DOWNTO 240) := ADC(11 DOWNTO 2);
			WHEN 25 => temp(259 DOWNTO 250) := ADC(11 DOWNTO 2);
			WHEN 26 => temp(269 DOWNTO 260) := ADC(11 DOWNTO 2);
			WHEN 27 => temp(279 DOWNTO 270) := ADC(11 DOWNTO 2);
			WHEN 28 => temp(289 DOWNTO 280) := ADC(11 DOWNTO 2);
			WHEN 29 => temp(299 DOWNTO 290) := ADC(11 DOWNTO 2);
			WHEN 30 => temp(309 DOWNTO 300) := ADC(11 DOWNTO 2);
			WHEN 31 => temp(319 DOWNTO 310) := ADC(11 DOWNTO 2);
			WHEN 32 => temp(329 DOWNTO 320) := ADC(11 DOWNTO 2);
			WHEN 33 => temp(339 DOWNTO 330) := ADC(11 DOWNTO 2);
			WHEN 34 => temp(349 DOWNTO 340) := ADC(11 DOWNTO 2);
			WHEN 35 => temp(359 DOWNTO 350) := ADC(11 DOWNTO 2);
			WHEN 36 => temp(369 DOWNTO 360) := ADC(11 DOWNTO 2);
			WHEN 37 => temp(379 DOWNTO 370) := ADC(11 DOWNTO 2);
			WHEN 38 => temp(389 DOWNTO 380) := ADC(11 DOWNTO 2);
			WHEN 39 => temp(399 DOWNTO 390) := ADC(11 DOWNTO 2);
			WHEN 40 => temp(409 DOWNTO 400) := ADC(11 DOWNTO 2);
			WHEN 41 => temp(419 DOWNTO 410) := ADC(11 DOWNTO 2);
			WHEN 42 => temp(429 DOWNTO 420) := ADC(11 DOWNTO 2);
			WHEN 43 => temp(439 DOWNTO 430) := ADC(11 DOWNTO 2);
			WHEN 44 => temp(449 DOWNTO 440) := ADC(11 DOWNTO 2);
			WHEN 45 => temp(459 DOWNTO 450) := ADC(11 DOWNTO 2);
			WHEN 46 => temp(469 DOWNTO 460) := ADC(11 DOWNTO 2);
			WHEN 47 => temp(479 DOWNTO 470) := ADC(11 DOWNTO 2);
			WHEN 48 => temp(489 DOWNTO 480) := ADC(11 DOWNTO 2);
			WHEN 49 => temp(499 DOWNTO 490) := ADC(11 DOWNTO 2);
			WHEN 50 => temp(509 DOWNTO 500) := ADC(11 DOWNTO 2);
			WHEN 51 => temp(519 DOWNTO 510) := ADC(11 DOWNTO 2);
			WHEN 52 => temp(529 DOWNTO 520) := ADC(11 DOWNTO 2);
			WHEN 53 => temp(539 DOWNTO 530) := ADC(11 DOWNTO 2);
			WHEN 54 => temp(549 DOWNTO 540) := ADC(11 DOWNTO 2);
			WHEN 55 => temp(559 DOWNTO 550) := ADC(11 DOWNTO 2);
			WHEN 56 => temp(569 DOWNTO 560) := ADC(11 DOWNTO 2);
			WHEN 57 => temp(579 DOWNTO 570) := ADC(11 DOWNTO 2);
			WHEN 58 => temp(589 DOWNTO 580) := ADC(11 DOWNTO 2);
			WHEN 59 => temp(599 DOWNTO 590) := ADC(11 DOWNTO 2);
			WHEN 60 => temp(609 DOWNTO 600) := ADC(11 DOWNTO 2);
			WHEN 61 => temp(619 DOWNTO 610) := ADC(11 DOWNTO 2);
			WHEN 62 => temp(629 DOWNTO 620) := ADC(11 DOWNTO 2);
			WHEN 63 => temp(639 DOWNTO 630) := ADC(11 DOWNTO 2);
			WHEN 64 => temp(649 DOWNTO 640) := ADC(11 DOWNTO 2);
			WHEN 65 => temp(659 DOWNTO 650) := ADC(11 DOWNTO 2);
			WHEN 66 => temp(669 DOWNTO 660) := ADC(11 DOWNTO 2);
			WHEN 67 => temp(679 DOWNTO 670) := ADC(11 DOWNTO 2);
			WHEN 68 => temp(689 DOWNTO 680) := ADC(11 DOWNTO 2);
			WHEN 69 => temp(699 DOWNTO 690) := ADC(11 DOWNTO 2);
			WHEN 70 => temp(709 DOWNTO 700) := ADC(11 DOWNTO 2);
			WHEN 71 => temp(719 DOWNTO 710) := ADC(11 DOWNTO 2);
			WHEN 72 => temp(729 DOWNTO 720) := ADC(11 DOWNTO 2);
			WHEN 73 => temp(739 DOWNTO 730) := ADC(11 DOWNTO 2);
			WHEN 74 => temp(749 DOWNTO 740) := ADC(11 DOWNTO 2);
			WHEN 75 => temp(759 DOWNTO 750) := ADC(11 DOWNTO 2);
			WHEN 76 => temp(769 DOWNTO 760) := ADC(11 DOWNTO 2);
			WHEN 77 => temp(779 DOWNTO 770) := ADC(11 DOWNTO 2);
			WHEN 78 => temp(789 DOWNTO 780) := ADC(11 DOWNTO 2);
			WHEN 79 => temp(799 DOWNTO 790) := ADC(11 DOWNTO 2);
			WHEN 80 => temp(809 DOWNTO 800) := ADC(11 DOWNTO 2);
			WHEN 81 => temp(819 DOWNTO 810) := ADC(11 DOWNTO 2);
			WHEN 82 => temp(829 DOWNTO 820) := ADC(11 DOWNTO 2);
			WHEN 83 => temp(839 DOWNTO 830) := ADC(11 DOWNTO 2);
			WHEN 84 => temp(849 DOWNTO 840) := ADC(11 DOWNTO 2);
			WHEN 85 => temp(859 DOWNTO 850) := ADC(11 DOWNTO 2);
			WHEN 86 => temp(869 DOWNTO 860) := ADC(11 DOWNTO 2);
			WHEN 87 => temp(879 DOWNTO 870) := ADC(11 DOWNTO 2);
			WHEN 88 => temp(889 DOWNTO 880) := ADC(11 DOWNTO 2);
			WHEN 89 => temp(899 DOWNTO 890) := ADC(11 DOWNTO 2);
			WHEN 90 => temp(909 DOWNTO 900) := ADC(11 DOWNTO 2);
			WHEN 91 => temp(919 DOWNTO 910) := ADC(11 DOWNTO 2);
			WHEN 92 => temp(929 DOWNTO 920) := ADC(11 DOWNTO 2);
			WHEN 93 => temp(939 DOWNTO 930) := ADC(11 DOWNTO 2);
			WHEN 94 => temp(949 DOWNTO 940) := ADC(11 DOWNTO 2);
			WHEN 95 => temp(959 DOWNTO 950) := ADC(11 DOWNTO 2);
			WHEN 96 => temp(969 DOWNTO 960) := ADC(11 DOWNTO 2);
			WHEN 97 => temp(979 DOWNTO 970) := ADC(11 DOWNTO 2);
			WHEN 98 => temp(989 DOWNTO 980) := ADC(11 DOWNTO 2);
			WHEN 99 => temp(999 DOWNTO 990) := ADC(11 DOWNTO 2);
			WHEN 100 => temp(1009 DOWNTO 1000) := ADC(11 DOWNTO 2);
			WHEN 101 => temp(1019 DOWNTO 1010) := ADC(11 DOWNTO 2);
			WHEN 102 => temp(1029 DOWNTO 1020) := ADC(11 DOWNTO 2);
			WHEN 103 => temp(1039 DOWNTO 1030) := ADC(11 DOWNTO 2);
			WHEN 104 => temp(1049 DOWNTO 1040) := ADC(11 DOWNTO 2);
			WHEN 105 => temp(1059 DOWNTO 1050) := ADC(11 DOWNTO 2);
			WHEN 106 => temp(1069 DOWNTO 1060) := ADC(11 DOWNTO 2);
			WHEN 107 => temp(1079 DOWNTO 1070) := ADC(11 DOWNTO 2);
			WHEN 108 => temp(1089 DOWNTO 1080) := ADC(11 DOWNTO 2);
			WHEN 109 => temp(1099 DOWNTO 1090) := ADC(11 DOWNTO 2);
			WHEN 110 => temp(1109 DOWNTO 1100) := ADC(11 DOWNTO 2);
			WHEN 111 => temp(1119 DOWNTO 1110) := ADC(11 DOWNTO 2);
			WHEN 112 => temp(1129 DOWNTO 1120) := ADC(11 DOWNTO 2);
			WHEN 113 => temp(1139 DOWNTO 1130) := ADC(11 DOWNTO 2);
			WHEN 114 => temp(1149 DOWNTO 1140) := ADC(11 DOWNTO 2);
			WHEN 115 => temp(1159 DOWNTO 1150) := ADC(11 DOWNTO 2);
			WHEN 116 => temp(1169 DOWNTO 1160) := ADC(11 DOWNTO 2);
			WHEN 117 => temp(1179 DOWNTO 1170) := ADC(11 DOWNTO 2);
			WHEN 118 => temp(1189 DOWNTO 1180) := ADC(11 DOWNTO 2);
			WHEN 119 => temp(1199 DOWNTO 1190) := ADC(11 DOWNTO 2);
			WHEN 120 => temp(1209 DOWNTO 1200) := ADC(11 DOWNTO 2);
			WHEN 121 => temp(1219 DOWNTO 1210) := ADC(11 DOWNTO 2);
			WHEN 122 => temp(1229 DOWNTO 1220) := ADC(11 DOWNTO 2);
			WHEN 123 => temp(1239 DOWNTO 1230) := ADC(11 DOWNTO 2);
			WHEN 124 => temp(1249 DOWNTO 1240) := ADC(11 DOWNTO 2);
			WHEN 125 => temp(1259 DOWNTO 1250) := ADC(11 DOWNTO 2);
			WHEN 126 => temp(1269 DOWNTO 1260) := ADC(11 DOWNTO 2);
			WHEN 127 => temp(1279 DOWNTO 1270) := ADC(11 DOWNTO 2);
			WHEN 128 => temp(1289 DOWNTO 1280) := ADC(11 DOWNTO 2);
			WHEN 129 => temp(1299 DOWNTO 1290) := ADC(11 DOWNTO 2);
			WHEN 130 => temp(1309 DOWNTO 1300) := ADC(11 DOWNTO 2);
			WHEN 131 => temp(1319 DOWNTO 1310) := ADC(11 DOWNTO 2);
			WHEN 132 => temp(1329 DOWNTO 1320) := ADC(11 DOWNTO 2);
			WHEN 133 => temp(1339 DOWNTO 1330) := ADC(11 DOWNTO 2);
			WHEN 134 => temp(1349 DOWNTO 1340) := ADC(11 DOWNTO 2);
			WHEN 135 => temp(1359 DOWNTO 1350) := ADC(11 DOWNTO 2);
			WHEN 136 => temp(1369 DOWNTO 1360) := ADC(11 DOWNTO 2);
			WHEN 137 => temp(1379 DOWNTO 1370) := ADC(11 DOWNTO 2);
			WHEN 138 => temp(1389 DOWNTO 1380) := ADC(11 DOWNTO 2);
			WHEN 139 => temp(1399 DOWNTO 1390) := ADC(11 DOWNTO 2);
			WHEN 140 => temp(1409 DOWNTO 1400) := ADC(11 DOWNTO 2);
			WHEN 141 => temp(1419 DOWNTO 1410) := ADC(11 DOWNTO 2);
			WHEN 142 => temp(1429 DOWNTO 1420) := ADC(11 DOWNTO 2);
			WHEN 143 => temp(1439 DOWNTO 1430) := ADC(11 DOWNTO 2);
			WHEN 144 => temp(1449 DOWNTO 1440) := ADC(11 DOWNTO 2);
			WHEN 145 => temp(1459 DOWNTO 1450) := ADC(11 DOWNTO 2);
			WHEN 146 => temp(1469 DOWNTO 1460) := ADC(11 DOWNTO 2);
			WHEN 147 => temp(1479 DOWNTO 1470) := ADC(11 DOWNTO 2);
			WHEN 148 => temp(1489 DOWNTO 1480) := ADC(11 DOWNTO 2);
			WHEN 149 => temp(1499 DOWNTO 1490) := ADC(11 DOWNTO 2);
			WHEN 150 => temp(1509 DOWNTO 1500) := ADC(11 DOWNTO 2);
			WHEN 151 => temp(1519 DOWNTO 1510) := ADC(11 DOWNTO 2);
			WHEN 152 => temp(1529 DOWNTO 1520) := ADC(11 DOWNTO 2);
			WHEN 153 => temp(1539 DOWNTO 1530) := ADC(11 DOWNTO 2);
			WHEN 154 => temp(1549 DOWNTO 1540) := ADC(11 DOWNTO 2);
			WHEN 155 => temp(1559 DOWNTO 1550) := ADC(11 DOWNTO 2);
			WHEN 156 => temp(1569 DOWNTO 1560) := ADC(11 DOWNTO 2);
			WHEN 157 => temp(1579 DOWNTO 1570) := ADC(11 DOWNTO 2);
			WHEN 158 => temp(1589 DOWNTO 1580) := ADC(11 DOWNTO 2);
			WHEN 159 => temp(1599 DOWNTO 1590) := ADC(11 DOWNTO 2);
			WHEN 160 => temp(1609 DOWNTO 1600) := ADC(11 DOWNTO 2);
			WHEN 161 => temp(1619 DOWNTO 1610) := ADC(11 DOWNTO 2);
			WHEN 162 => temp(1629 DOWNTO 1620) := ADC(11 DOWNTO 2);
			WHEN 163 => temp(1639 DOWNTO 1630) := ADC(11 DOWNTO 2);
			WHEN 164 => temp(1649 DOWNTO 1640) := ADC(11 DOWNTO 2);
			WHEN 165 => temp(1659 DOWNTO 1650) := ADC(11 DOWNTO 2);
			WHEN 166 => temp(1669 DOWNTO 1660) := ADC(11 DOWNTO 2);
			WHEN 167 => temp(1679 DOWNTO 1670) := ADC(11 DOWNTO 2);
			WHEN 168 => temp(1689 DOWNTO 1680) := ADC(11 DOWNTO 2);
			WHEN 169 => temp(1699 DOWNTO 1690) := ADC(11 DOWNTO 2);
			WHEN 170 => temp(1709 DOWNTO 1700) := ADC(11 DOWNTO 2);
			WHEN 171 => temp(1719 DOWNTO 1710) := ADC(11 DOWNTO 2);
			WHEN 172 => temp(1729 DOWNTO 1720) := ADC(11 DOWNTO 2);
			WHEN 173 => temp(1739 DOWNTO 1730) := ADC(11 DOWNTO 2);
			WHEN 174 => temp(1749 DOWNTO 1740) := ADC(11 DOWNTO 2);
			WHEN 175 => temp(1759 DOWNTO 1750) := ADC(11 DOWNTO 2);
			WHEN 176 => temp(1769 DOWNTO 1760) := ADC(11 DOWNTO 2);
			WHEN 177 => temp(1779 DOWNTO 1770) := ADC(11 DOWNTO 2);
			WHEN 178 => temp(1789 DOWNTO 1780) := ADC(11 DOWNTO 2);
			WHEN 179 => temp(1799 DOWNTO 1790) := ADC(11 DOWNTO 2);
			WHEN 180 => temp(1809 DOWNTO 1800) := ADC(11 DOWNTO 2);
			WHEN 181 => temp(1819 DOWNTO 1810) := ADC(11 DOWNTO 2);
			WHEN 182 => temp(1829 DOWNTO 1820) := ADC(11 DOWNTO 2);
			WHEN 183 => temp(1839 DOWNTO 1830) := ADC(11 DOWNTO 2);
			WHEN 184 => temp(1849 DOWNTO 1840) := ADC(11 DOWNTO 2);
			WHEN 185 => temp(1859 DOWNTO 1850) := ADC(11 DOWNTO 2);
			WHEN 186 => temp(1869 DOWNTO 1860) := ADC(11 DOWNTO 2);
			WHEN 187 => temp(1879 DOWNTO 1870) := ADC(11 DOWNTO 2);
			WHEN 188 => temp(1889 DOWNTO 1880) := ADC(11 DOWNTO 2);
			WHEN 189 => temp(1899 DOWNTO 1890) := ADC(11 DOWNTO 2);
			WHEN 190 => temp(1909 DOWNTO 1900) := ADC(11 DOWNTO 2);
			WHEN 191 => temp(1919 DOWNTO 1910) := ADC(11 DOWNTO 2);
			WHEN 192 => temp(1929 DOWNTO 1920) := ADC(11 DOWNTO 2);
			WHEN 193 => temp(1939 DOWNTO 1930) := ADC(11 DOWNTO 2);
			WHEN 194 => temp(1949 DOWNTO 1940) := ADC(11 DOWNTO 2);
			WHEN 195 => temp(1959 DOWNTO 1950) := ADC(11 DOWNTO 2);
			WHEN 196 => temp(1969 DOWNTO 1960) := ADC(11 DOWNTO 2);
			WHEN 197 => temp(1979 DOWNTO 1970) := ADC(11 DOWNTO 2);
			WHEN 198 => temp(1989 DOWNTO 1980) := ADC(11 DOWNTO 2);
			WHEN 199 => temp(1999 DOWNTO 1990) := ADC(11 DOWNTO 2);
			WHEN 200 => temp(2009 DOWNTO 2000) := ADC(11 DOWNTO 2);
			WHEN 201 => temp(2019 DOWNTO 2010) := ADC(11 DOWNTO 2);
			WHEN 202 => temp(2029 DOWNTO 2020) := ADC(11 DOWNTO 2);
			WHEN 203 => temp(2039 DOWNTO 2030) := ADC(11 DOWNTO 2);
			WHEN 204 => temp(2049 DOWNTO 2040) := ADC(11 DOWNTO 2);
			WHEN 205 => temp(2059 DOWNTO 2050) := ADC(11 DOWNTO 2);
			WHEN 206 => temp(2069 DOWNTO 2060) := ADC(11 DOWNTO 2);
			WHEN 207 => temp(2079 DOWNTO 2070) := ADC(11 DOWNTO 2);
			WHEN 208 => temp(2089 DOWNTO 2080) := ADC(11 DOWNTO 2);
			WHEN 209 => temp(2099 DOWNTO 2090) := ADC(11 DOWNTO 2);
			WHEN 210 => temp(2109 DOWNTO 2100) := ADC(11 DOWNTO 2);
			WHEN 211 => temp(2119 DOWNTO 2110) := ADC(11 DOWNTO 2);
			WHEN 212 => temp(2129 DOWNTO 2120) := ADC(11 DOWNTO 2);
			WHEN 213 => temp(2139 DOWNTO 2130) := ADC(11 DOWNTO 2);
			WHEN 214 => temp(2149 DOWNTO 2140) := ADC(11 DOWNTO 2);
			WHEN 215 => temp(2159 DOWNTO 2150) := ADC(11 DOWNTO 2);
			WHEN 216 => temp(2169 DOWNTO 2160) := ADC(11 DOWNTO 2);
			WHEN 217 => temp(2179 DOWNTO 2170) := ADC(11 DOWNTO 2);
			WHEN 218 => temp(2189 DOWNTO 2180) := ADC(11 DOWNTO 2);
			WHEN 219 => temp(2199 DOWNTO 2190) := ADC(11 DOWNTO 2);
			WHEN 220 => temp(2209 DOWNTO 2200) := ADC(11 DOWNTO 2);
			WHEN 221 => temp(2219 DOWNTO 2210) := ADC(11 DOWNTO 2);
			WHEN 222 => temp(2229 DOWNTO 2220) := ADC(11 DOWNTO 2);
			WHEN 223 => temp(2239 DOWNTO 2230) := ADC(11 DOWNTO 2);
			WHEN 224 => temp(2249 DOWNTO 2240) := ADC(11 DOWNTO 2);
			WHEN 225 => temp(2259 DOWNTO 2250) := ADC(11 DOWNTO 2);
			WHEN 226 => temp(2269 DOWNTO 2260) := ADC(11 DOWNTO 2);
			WHEN 227 => temp(2279 DOWNTO 2270) := ADC(11 DOWNTO 2);
			WHEN 228 => temp(2289 DOWNTO 2280) := ADC(11 DOWNTO 2);
			WHEN 229 => temp(2299 DOWNTO 2290) := ADC(11 DOWNTO 2);
			WHEN 230 => temp(2309 DOWNTO 2300) := ADC(11 DOWNTO 2);
			WHEN 231 => temp(2319 DOWNTO 2310) := ADC(11 DOWNTO 2);
			WHEN 232 => temp(2329 DOWNTO 2320) := ADC(11 DOWNTO 2);
			WHEN 233 => temp(2339 DOWNTO 2330) := ADC(11 DOWNTO 2);
			WHEN 234 => temp(2349 DOWNTO 2340) := ADC(11 DOWNTO 2);
			WHEN 235 => temp(2359 DOWNTO 2350) := ADC(11 DOWNTO 2);
			WHEN 236 => temp(2369 DOWNTO 2360) := ADC(11 DOWNTO 2);
			WHEN 237 => temp(2379 DOWNTO 2370) := ADC(11 DOWNTO 2);
			WHEN 238 => temp(2389 DOWNTO 2380) := ADC(11 DOWNTO 2);
			WHEN 239 => temp(2399 DOWNTO 2390) := ADC(11 DOWNTO 2);
			WHEN 240 => temp(2409 DOWNTO 2400) := ADC(11 DOWNTO 2);
			WHEN 241 => temp(2419 DOWNTO 2410) := ADC(11 DOWNTO 2);
			WHEN 242 => temp(2429 DOWNTO 2420) := ADC(11 DOWNTO 2);
			WHEN 243 => temp(2439 DOWNTO 2430) := ADC(11 DOWNTO 2);
			WHEN 244 => temp(2449 DOWNTO 2440) := ADC(11 DOWNTO 2);
			WHEN 245 => temp(2459 DOWNTO 2450) := ADC(11 DOWNTO 2);
			WHEN 246 => temp(2469 DOWNTO 2460) := ADC(11 DOWNTO 2);
			WHEN 247 => temp(2479 DOWNTO 2470) := ADC(11 DOWNTO 2);
			WHEN 248 => temp(2489 DOWNTO 2480) := ADC(11 DOWNTO 2);
			WHEN 249 => temp(2499 DOWNTO 2490) := ADC(11 DOWNTO 2);
			WHEN 250 => temp(2509 DOWNTO 2500) := ADC(11 DOWNTO 2);
			WHEN 251 => temp(2519 DOWNTO 2510) := ADC(11 DOWNTO 2);
			WHEN 252 => temp(2529 DOWNTO 2520) := ADC(11 DOWNTO 2);
			WHEN 253 => temp(2539 DOWNTO 2530) := ADC(11 DOWNTO 2);
			WHEN 254 => temp(2549 DOWNTO 2540) := ADC(11 DOWNTO 2);
			WHEN 255 => temp(2559 DOWNTO 2550) := ADC(11 DOWNTO 2);
			WHEN 256 => temp(2569 DOWNTO 2560) := ADC(11 DOWNTO 2);
			WHEN 257 => temp(2579 DOWNTO 2570) := ADC(11 DOWNTO 2);
			WHEN 258 => temp(2589 DOWNTO 2580) := ADC(11 DOWNTO 2);
			WHEN 259 => temp(2599 DOWNTO 2590) := ADC(11 DOWNTO 2);
			WHEN 260 => temp(2609 DOWNTO 2600) := ADC(11 DOWNTO 2);
			WHEN 261 => temp(2619 DOWNTO 2610) := ADC(11 DOWNTO 2);
			WHEN 262 => temp(2629 DOWNTO 2620) := ADC(11 DOWNTO 2);
			WHEN 263 => temp(2639 DOWNTO 2630) := ADC(11 DOWNTO 2);
			WHEN 264 => temp(2649 DOWNTO 2640) := ADC(11 DOWNTO 2);
			WHEN 265 => temp(2659 DOWNTO 2650) := ADC(11 DOWNTO 2);
			WHEN 266 => temp(2669 DOWNTO 2660) := ADC(11 DOWNTO 2);
			WHEN 267 => temp(2679 DOWNTO 2670) := ADC(11 DOWNTO 2);
			WHEN 268 => temp(2689 DOWNTO 2680) := ADC(11 DOWNTO 2);
			WHEN 269 => temp(2699 DOWNTO 2690) := ADC(11 DOWNTO 2);
			WHEN 270 => temp(2709 DOWNTO 2700) := ADC(11 DOWNTO 2);
			WHEN 271 => temp(2719 DOWNTO 2710) := ADC(11 DOWNTO 2);
			WHEN 272 => temp(2729 DOWNTO 2720) := ADC(11 DOWNTO 2);
			WHEN 273 => temp(2739 DOWNTO 2730) := ADC(11 DOWNTO 2);
			WHEN 274 => temp(2749 DOWNTO 2740) := ADC(11 DOWNTO 2);
			WHEN 275 => temp(2759 DOWNTO 2750) := ADC(11 DOWNTO 2);
			WHEN 276 => temp(2769 DOWNTO 2760) := ADC(11 DOWNTO 2);
			WHEN 277 => temp(2779 DOWNTO 2770) := ADC(11 DOWNTO 2);
			WHEN 278 => temp(2789 DOWNTO 2780) := ADC(11 DOWNTO 2);
			WHEN 279 => temp(2799 DOWNTO 2790) := ADC(11 DOWNTO 2);
			WHEN 280 => temp(2809 DOWNTO 2800) := ADC(11 DOWNTO 2);
			WHEN 281 => temp(2819 DOWNTO 2810) := ADC(11 DOWNTO 2);
			WHEN 282 => temp(2829 DOWNTO 2820) := ADC(11 DOWNTO 2);
			WHEN 283 => temp(2839 DOWNTO 2830) := ADC(11 DOWNTO 2);
			WHEN 284 => temp(2849 DOWNTO 2840) := ADC(11 DOWNTO 2);
			WHEN 285 => temp(2859 DOWNTO 2850) := ADC(11 DOWNTO 2);
			WHEN 286 => temp(2869 DOWNTO 2860) := ADC(11 DOWNTO 2);
			WHEN 287 => temp(2879 DOWNTO 2870) := ADC(11 DOWNTO 2);
			WHEN 288 => temp(2889 DOWNTO 2880) := ADC(11 DOWNTO 2);
			WHEN 289 => temp(2899 DOWNTO 2890) := ADC(11 DOWNTO 2);
			WHEN 290 => temp(2909 DOWNTO 2900) := ADC(11 DOWNTO 2);
			WHEN 291 => temp(2919 DOWNTO 2910) := ADC(11 DOWNTO 2);
			WHEN 292 => temp(2929 DOWNTO 2920) := ADC(11 DOWNTO 2);
			WHEN 293 => temp(2939 DOWNTO 2930) := ADC(11 DOWNTO 2);
			WHEN 294 => temp(2949 DOWNTO 2940) := ADC(11 DOWNTO 2);
			WHEN 295 => temp(2959 DOWNTO 2950) := ADC(11 DOWNTO 2);
			WHEN 296 => temp(2969 DOWNTO 2960) := ADC(11 DOWNTO 2);
			WHEN 297 => temp(2979 DOWNTO 2970) := ADC(11 DOWNTO 2);
			WHEN 298 => temp(2989 DOWNTO 2980) := ADC(11 DOWNTO 2);
			WHEN 299 => temp(2999 DOWNTO 2990) := ADC(11 DOWNTO 2);
			WHEN 300 => temp(3009 DOWNTO 3000) := ADC(11 DOWNTO 2);
			WHEN 301 => temp(3019 DOWNTO 3010) := ADC(11 DOWNTO 2);
			WHEN 302 => temp(3029 DOWNTO 3020) := ADC(11 DOWNTO 2);
			WHEN 303 => temp(3039 DOWNTO 3030) := ADC(11 DOWNTO 2);
			WHEN 304 => temp(3049 DOWNTO 3040) := ADC(11 DOWNTO 2);
			WHEN 305 => temp(3059 DOWNTO 3050) := ADC(11 DOWNTO 2);
			WHEN 306 => temp(3069 DOWNTO 3060) := ADC(11 DOWNTO 2);
			WHEN 307 => temp(3079 DOWNTO 3070) := ADC(11 DOWNTO 2);
			WHEN 308 => temp(3089 DOWNTO 3080) := ADC(11 DOWNTO 2);
			WHEN 309 => temp(3099 DOWNTO 3090) := ADC(11 DOWNTO 2);
			WHEN 310 => temp(3109 DOWNTO 3100) := ADC(11 DOWNTO 2);
			WHEN 311 => temp(3119 DOWNTO 3110) := ADC(11 DOWNTO 2);
			WHEN 312 => temp(3129 DOWNTO 3120) := ADC(11 DOWNTO 2);
			WHEN 313 => temp(3139 DOWNTO 3130) := ADC(11 DOWNTO 2);
			WHEN 314 => temp(3149 DOWNTO 3140) := ADC(11 DOWNTO 2);
			WHEN 315 => temp(3159 DOWNTO 3150) := ADC(11 DOWNTO 2);
			WHEN 316 => temp(3169 DOWNTO 3160) := ADC(11 DOWNTO 2);
			WHEN 317 => temp(3179 DOWNTO 3170) := ADC(11 DOWNTO 2);
			WHEN 318 => temp(3189 DOWNTO 3180) := ADC(11 DOWNTO 2);
			WHEN 319 => temp(3199 DOWNTO 3190) := ADC(11 DOWNTO 2);
			WHEN 320 => temp(3209 DOWNTO 3200) := ADC(11 DOWNTO 2);
			WHEN 321 => temp(3219 DOWNTO 3210) := ADC(11 DOWNTO 2);
			WHEN 322 => temp(3229 DOWNTO 3220) := ADC(11 DOWNTO 2);
			WHEN 323 => temp(3239 DOWNTO 3230) := ADC(11 DOWNTO 2);
			WHEN 324 => temp(3249 DOWNTO 3240) := ADC(11 DOWNTO 2);
			WHEN 325 => temp(3259 DOWNTO 3250) := ADC(11 DOWNTO 2);
			WHEN 326 => temp(3269 DOWNTO 3260) := ADC(11 DOWNTO 2);
			WHEN 327 => temp(3279 DOWNTO 3270) := ADC(11 DOWNTO 2);
			WHEN 328 => temp(3289 DOWNTO 3280) := ADC(11 DOWNTO 2);
			WHEN 329 => temp(3299 DOWNTO 3290) := ADC(11 DOWNTO 2);
			WHEN 330 => temp(3309 DOWNTO 3300) := ADC(11 DOWNTO 2);
			WHEN 331 => temp(3319 DOWNTO 3310) := ADC(11 DOWNTO 2);
			WHEN 332 => temp(3329 DOWNTO 3320) := ADC(11 DOWNTO 2);
			WHEN 333 => temp(3339 DOWNTO 3330) := ADC(11 DOWNTO 2);
			WHEN 334 => temp(3349 DOWNTO 3340) := ADC(11 DOWNTO 2);
			WHEN 335 => temp(3359 DOWNTO 3350) := ADC(11 DOWNTO 2);
			WHEN 336 => temp(3369 DOWNTO 3360) := ADC(11 DOWNTO 2);
			WHEN 337 => temp(3379 DOWNTO 3370) := ADC(11 DOWNTO 2);
			WHEN 338 => temp(3389 DOWNTO 3380) := ADC(11 DOWNTO 2);
			WHEN 339 => temp(3399 DOWNTO 3390) := ADC(11 DOWNTO 2);
			WHEN 340 => temp(3409 DOWNTO 3400) := ADC(11 DOWNTO 2);
			WHEN 341 => temp(3419 DOWNTO 3410) := ADC(11 DOWNTO 2);
			WHEN 342 => temp(3429 DOWNTO 3420) := ADC(11 DOWNTO 2);
			WHEN 343 => temp(3439 DOWNTO 3430) := ADC(11 DOWNTO 2);
			WHEN 344 => temp(3449 DOWNTO 3440) := ADC(11 DOWNTO 2);
			WHEN 345 => temp(3459 DOWNTO 3450) := ADC(11 DOWNTO 2);
			WHEN 346 => temp(3469 DOWNTO 3460) := ADC(11 DOWNTO 2);
			WHEN 347 => temp(3479 DOWNTO 3470) := ADC(11 DOWNTO 2);
			WHEN 348 => temp(3489 DOWNTO 3480) := ADC(11 DOWNTO 2);
			WHEN 349 => temp(3499 DOWNTO 3490) := ADC(11 DOWNTO 2);
			WHEN 350 => temp(3509 DOWNTO 3500) := ADC(11 DOWNTO 2);
			WHEN 351 => temp(3519 DOWNTO 3510) := ADC(11 DOWNTO 2);
			WHEN 352 => temp(3529 DOWNTO 3520) := ADC(11 DOWNTO 2);
			WHEN 353 => temp(3539 DOWNTO 3530) := ADC(11 DOWNTO 2);
			WHEN 354 => temp(3549 DOWNTO 3540) := ADC(11 DOWNTO 2);
			WHEN 355 => temp(3559 DOWNTO 3550) := ADC(11 DOWNTO 2);
			WHEN 356 => temp(3569 DOWNTO 3560) := ADC(11 DOWNTO 2);
			WHEN 357 => temp(3579 DOWNTO 3570) := ADC(11 DOWNTO 2);
			WHEN 358 => temp(3589 DOWNTO 3580) := ADC(11 DOWNTO 2);
			WHEN 359 => temp(3599 DOWNTO 3590) := ADC(11 DOWNTO 2);
			WHEN 360 => temp(3609 DOWNTO 3600) := ADC(11 DOWNTO 2);
			WHEN 361 => temp(3619 DOWNTO 3610) := ADC(11 DOWNTO 2);
			WHEN 362 => temp(3629 DOWNTO 3620) := ADC(11 DOWNTO 2);
			WHEN 363 => temp(3639 DOWNTO 3630) := ADC(11 DOWNTO 2);
			WHEN 364 => temp(3649 DOWNTO 3640) := ADC(11 DOWNTO 2);
			WHEN 365 => temp(3659 DOWNTO 3650) := ADC(11 DOWNTO 2);
			WHEN 366 => temp(3669 DOWNTO 3660) := ADC(11 DOWNTO 2);
			WHEN 367 => temp(3679 DOWNTO 3670) := ADC(11 DOWNTO 2);
			WHEN 368 => temp(3689 DOWNTO 3680) := ADC(11 DOWNTO 2);
			WHEN 369 => temp(3699 DOWNTO 3690) := ADC(11 DOWNTO 2);
			WHEN 370 => temp(3709 DOWNTO 3700) := ADC(11 DOWNTO 2);
			WHEN 371 => temp(3719 DOWNTO 3710) := ADC(11 DOWNTO 2);
			WHEN 372 => temp(3729 DOWNTO 3720) := ADC(11 DOWNTO 2);
			WHEN 373 => temp(3739 DOWNTO 3730) := ADC(11 DOWNTO 2);
			WHEN 374 => temp(3749 DOWNTO 3740) := ADC(11 DOWNTO 2);
			WHEN 375 => temp(3759 DOWNTO 3750) := ADC(11 DOWNTO 2);
			WHEN 376 => temp(3769 DOWNTO 3760) := ADC(11 DOWNTO 2);
			WHEN 377 => temp(3779 DOWNTO 3770) := ADC(11 DOWNTO 2);
			WHEN 378 => temp(3789 DOWNTO 3780) := ADC(11 DOWNTO 2);
			WHEN 379 => temp(3799 DOWNTO 3790) := ADC(11 DOWNTO 2);
			WHEN 380 => temp(3809 DOWNTO 3800) := ADC(11 DOWNTO 2);
			WHEN 381 => temp(3819 DOWNTO 3810) := ADC(11 DOWNTO 2);
			WHEN 382 => temp(3829 DOWNTO 3820) := ADC(11 DOWNTO 2);
			WHEN 383 => temp(3839 DOWNTO 3830) := ADC(11 DOWNTO 2);
			WHEN 384 => temp(3849 DOWNTO 3840) := ADC(11 DOWNTO 2);
			WHEN 385 => temp(3859 DOWNTO 3850) := ADC(11 DOWNTO 2);
			WHEN 386 => temp(3869 DOWNTO 3860) := ADC(11 DOWNTO 2);
			WHEN 387 => temp(3879 DOWNTO 3870) := ADC(11 DOWNTO 2);
			WHEN 388 => temp(3889 DOWNTO 3880) := ADC(11 DOWNTO 2);
			WHEN 389 => temp(3899 DOWNTO 3890) := ADC(11 DOWNTO 2);
			WHEN 390 => temp(3909 DOWNTO 3900) := ADC(11 DOWNTO 2);
			WHEN 391 => temp(3919 DOWNTO 3910) := ADC(11 DOWNTO 2);
			WHEN 392 => temp(3929 DOWNTO 3920) := ADC(11 DOWNTO 2);
			WHEN 393 => temp(3939 DOWNTO 3930) := ADC(11 DOWNTO 2);
			WHEN 394 => temp(3949 DOWNTO 3940) := ADC(11 DOWNTO 2);
			WHEN 395 => temp(3959 DOWNTO 3950) := ADC(11 DOWNTO 2);
			WHEN 396 => temp(3969 DOWNTO 3960) := ADC(11 DOWNTO 2);
			WHEN 397 => temp(3979 DOWNTO 3970) := ADC(11 DOWNTO 2);
			WHEN 398 => temp(3989 DOWNTO 3980) := ADC(11 DOWNTO 2);
			WHEN 399 => temp(3999 DOWNTO 3990) := ADC(11 DOWNTO 2);
			WHEN 400 => temp(4009 DOWNTO 4000) := ADC(11 DOWNTO 2);
			WHEN 401 => temp(4019 DOWNTO 4010) := ADC(11 DOWNTO 2);
			WHEN 402 => temp(4029 DOWNTO 4020) := ADC(11 DOWNTO 2);
			WHEN 403 => temp(4039 DOWNTO 4030) := ADC(11 DOWNTO 2);
			WHEN 404 => temp(4049 DOWNTO 4040) := ADC(11 DOWNTO 2);
			WHEN 405 => temp(4059 DOWNTO 4050) := ADC(11 DOWNTO 2);
			WHEN 406 => temp(4069 DOWNTO 4060) := ADC(11 DOWNTO 2);
			WHEN 407 => temp(4079 DOWNTO 4070) := ADC(11 DOWNTO 2);
			WHEN 408 => temp(4089 DOWNTO 4080) := ADC(11 DOWNTO 2);
			WHEN 409 => temp(4099 DOWNTO 4090) := ADC(11 DOWNTO 2);
			WHEN 410 => temp(4109 DOWNTO 4100) := ADC(11 DOWNTO 2);
			WHEN 411 => temp(4119 DOWNTO 4110) := ADC(11 DOWNTO 2);
			WHEN 412 => temp(4129 DOWNTO 4120) := ADC(11 DOWNTO 2);
			WHEN 413 => temp(4139 DOWNTO 4130) := ADC(11 DOWNTO 2);
			WHEN 414 => temp(4149 DOWNTO 4140) := ADC(11 DOWNTO 2);
			WHEN 415 => temp(4159 DOWNTO 4150) := ADC(11 DOWNTO 2);
			WHEN 416 => temp(4169 DOWNTO 4160) := ADC(11 DOWNTO 2);
			WHEN 417 => temp(4179 DOWNTO 4170) := ADC(11 DOWNTO 2);
			WHEN 418 => temp(4189 DOWNTO 4180) := ADC(11 DOWNTO 2);
			WHEN 419 => temp(4199 DOWNTO 4190) := ADC(11 DOWNTO 2);
			WHEN 420 => temp(4209 DOWNTO 4200) := ADC(11 DOWNTO 2);
			WHEN 421 => temp(4219 DOWNTO 4210) := ADC(11 DOWNTO 2);
			WHEN 422 => temp(4229 DOWNTO 4220) := ADC(11 DOWNTO 2);
			WHEN 423 => temp(4239 DOWNTO 4230) := ADC(11 DOWNTO 2);
			WHEN 424 => temp(4249 DOWNTO 4240) := ADC(11 DOWNTO 2);
			WHEN 425 => temp(4259 DOWNTO 4250) := ADC(11 DOWNTO 2);
			WHEN 426 => temp(4269 DOWNTO 4260) := ADC(11 DOWNTO 2);
			WHEN 427 => temp(4279 DOWNTO 4270) := ADC(11 DOWNTO 2);
			WHEN 428 => temp(4289 DOWNTO 4280) := ADC(11 DOWNTO 2);
			WHEN 429 => temp(4299 DOWNTO 4290) := ADC(11 DOWNTO 2);
			WHEN 430 => temp(4309 DOWNTO 4300) := ADC(11 DOWNTO 2);
			WHEN 431 => temp(4319 DOWNTO 4310) := ADC(11 DOWNTO 2);
			WHEN 432 => temp(4329 DOWNTO 4320) := ADC(11 DOWNTO 2);
			WHEN 433 => temp(4339 DOWNTO 4330) := ADC(11 DOWNTO 2);
			WHEN 434 => temp(4349 DOWNTO 4340) := ADC(11 DOWNTO 2);
			WHEN 435 => temp(4359 DOWNTO 4350) := ADC(11 DOWNTO 2);
			WHEN 436 => temp(4369 DOWNTO 4360) := ADC(11 DOWNTO 2);
			WHEN 437 => temp(4379 DOWNTO 4370) := ADC(11 DOWNTO 2);
			WHEN 438 => temp(4389 DOWNTO 4380) := ADC(11 DOWNTO 2);
			WHEN 439 => temp(4399 DOWNTO 4390) := ADC(11 DOWNTO 2);
			WHEN 440 => temp(4409 DOWNTO 4400) := ADC(11 DOWNTO 2);
			WHEN 441 => temp(4419 DOWNTO 4410) := ADC(11 DOWNTO 2);
			WHEN 442 => temp(4429 DOWNTO 4420) := ADC(11 DOWNTO 2);
			WHEN 443 => temp(4439 DOWNTO 4430) := ADC(11 DOWNTO 2);
			WHEN 444 => temp(4449 DOWNTO 4440) := ADC(11 DOWNTO 2);
			WHEN 445 => temp(4459 DOWNTO 4450) := ADC(11 DOWNTO 2);
			WHEN 446 => temp(4469 DOWNTO 4460) := ADC(11 DOWNTO 2);
			WHEN 447 => temp(4479 DOWNTO 4470) := ADC(11 DOWNTO 2);
			WHEN 448 => temp(4489 DOWNTO 4480) := ADC(11 DOWNTO 2);
			WHEN 449 => temp(4499 DOWNTO 4490) := ADC(11 DOWNTO 2);
			WHEN 450 => temp(4509 DOWNTO 4500) := ADC(11 DOWNTO 2);
			WHEN 451 => temp(4519 DOWNTO 4510) := ADC(11 DOWNTO 2);
			WHEN 452 => temp(4529 DOWNTO 4520) := ADC(11 DOWNTO 2);
			WHEN 453 => temp(4539 DOWNTO 4530) := ADC(11 DOWNTO 2);
			WHEN 454 => temp(4549 DOWNTO 4540) := ADC(11 DOWNTO 2);
			WHEN 455 => temp(4559 DOWNTO 4550) := ADC(11 DOWNTO 2);
			WHEN 456 => temp(4569 DOWNTO 4560) := ADC(11 DOWNTO 2);
			WHEN 457 => temp(4579 DOWNTO 4570) := ADC(11 DOWNTO 2);
			WHEN 458 => temp(4589 DOWNTO 4580) := ADC(11 DOWNTO 2);
			WHEN 459 => temp(4599 DOWNTO 4590) := ADC(11 DOWNTO 2);
			WHEN 460 => temp(4609 DOWNTO 4600) := ADC(11 DOWNTO 2);
			WHEN 461 => temp(4619 DOWNTO 4610) := ADC(11 DOWNTO 2);
			WHEN 462 => temp(4629 DOWNTO 4620) := ADC(11 DOWNTO 2);
			WHEN 463 => temp(4639 DOWNTO 4630) := ADC(11 DOWNTO 2);
			WHEN 464 => temp(4649 DOWNTO 4640) := ADC(11 DOWNTO 2);
			WHEN 465 => temp(4659 DOWNTO 4650) := ADC(11 DOWNTO 2);
			WHEN 466 => temp(4669 DOWNTO 4660) := ADC(11 DOWNTO 2);
			WHEN 467 => temp(4679 DOWNTO 4670) := ADC(11 DOWNTO 2);
			WHEN 468 => temp(4689 DOWNTO 4680) := ADC(11 DOWNTO 2);
			WHEN 469 => temp(4699 DOWNTO 4690) := ADC(11 DOWNTO 2);
			WHEN 470 => temp(4709 DOWNTO 4700) := ADC(11 DOWNTO 2);
			WHEN 471 => temp(4719 DOWNTO 4710) := ADC(11 DOWNTO 2);
			WHEN 472 => temp(4729 DOWNTO 4720) := ADC(11 DOWNTO 2);
			WHEN 473 => temp(4739 DOWNTO 4730) := ADC(11 DOWNTO 2);
			WHEN 474 => temp(4749 DOWNTO 4740) := ADC(11 DOWNTO 2);
			WHEN 475 => temp(4759 DOWNTO 4750) := ADC(11 DOWNTO 2);
			WHEN 476 => temp(4769 DOWNTO 4760) := ADC(11 DOWNTO 2);
			WHEN 477 => temp(4779 DOWNTO 4770) := ADC(11 DOWNTO 2);
			WHEN 478 => temp(4789 DOWNTO 4780) := ADC(11 DOWNTO 2);
			WHEN 479 => temp(4799 DOWNTO 4790) := ADC(11 DOWNTO 2);
			WHEN 480 => temp(4809 DOWNTO 4800) := ADC(11 DOWNTO 2);
			WHEN 481 => temp(4819 DOWNTO 4810) := ADC(11 DOWNTO 2);
			WHEN 482 => temp(4829 DOWNTO 4820) := ADC(11 DOWNTO 2);
			WHEN 483 => temp(4839 DOWNTO 4830) := ADC(11 DOWNTO 2);
			WHEN 484 => temp(4849 DOWNTO 4840) := ADC(11 DOWNTO 2);
			WHEN 485 => temp(4859 DOWNTO 4850) := ADC(11 DOWNTO 2);
			WHEN 486 => temp(4869 DOWNTO 4860) := ADC(11 DOWNTO 2);
			WHEN 487 => temp(4879 DOWNTO 4870) := ADC(11 DOWNTO 2);
			WHEN 488 => temp(4889 DOWNTO 4880) := ADC(11 DOWNTO 2);
			WHEN 489 => temp(4899 DOWNTO 4890) := ADC(11 DOWNTO 2);
			WHEN 490 => temp(4909 DOWNTO 4900) := ADC(11 DOWNTO 2);
			WHEN 491 => temp(4919 DOWNTO 4910) := ADC(11 DOWNTO 2);
			WHEN 492 => temp(4929 DOWNTO 4920) := ADC(11 DOWNTO 2);
			WHEN 493 => temp(4939 DOWNTO 4930) := ADC(11 DOWNTO 2);
			WHEN 494 => temp(4949 DOWNTO 4940) := ADC(11 DOWNTO 2);
			WHEN 495 => temp(4959 DOWNTO 4950) := ADC(11 DOWNTO 2);
			WHEN 496 => temp(4969 DOWNTO 4960) := ADC(11 DOWNTO 2);
			WHEN 497 => temp(4979 DOWNTO 4970) := ADC(11 DOWNTO 2);
			WHEN 498 => temp(4989 DOWNTO 4980) := ADC(11 DOWNTO 2);
			WHEN 499 => temp(4999 DOWNTO 4990) := ADC(11 DOWNTO 2);
			WHEN 500 => temp(5009 DOWNTO 5000) := ADC(11 DOWNTO 2);
			WHEN 501 => temp(5019 DOWNTO 5010) := ADC(11 DOWNTO 2);
			WHEN 502 => temp(5029 DOWNTO 5020) := ADC(11 DOWNTO 2);
			WHEN 503 => temp(5039 DOWNTO 5030) := ADC(11 DOWNTO 2);
			WHEN 504 => temp(5049 DOWNTO 5040) := ADC(11 DOWNTO 2);
			WHEN 505 => temp(5059 DOWNTO 5050) := ADC(11 DOWNTO 2);
			WHEN 506 => temp(5069 DOWNTO 5060) := ADC(11 DOWNTO 2);
			WHEN 507 => temp(5079 DOWNTO 5070) := ADC(11 DOWNTO 2);
			WHEN 508 => temp(5089 DOWNTO 5080) := ADC(11 DOWNTO 2);
			WHEN 509 => temp(5099 DOWNTO 5090) := ADC(11 DOWNTO 2);
			WHEN 510 => temp(5109 DOWNTO 5100) := ADC(11 DOWNTO 2);
			WHEN 511 => temp(5119 DOWNTO 5110) := ADC(11 DOWNTO 2);
			WHEN 512 => temp(5129 DOWNTO 5120) := ADC(11 DOWNTO 2);
			WHEN 513 => temp(5139 DOWNTO 5130) := ADC(11 DOWNTO 2);
			WHEN 514 => temp(5149 DOWNTO 5140) := ADC(11 DOWNTO 2);
			WHEN 515 => temp(5159 DOWNTO 5150) := ADC(11 DOWNTO 2);
			WHEN 516 => temp(5169 DOWNTO 5160) := ADC(11 DOWNTO 2);
			WHEN 517 => temp(5179 DOWNTO 5170) := ADC(11 DOWNTO 2);
			WHEN 518 => temp(5189 DOWNTO 5180) := ADC(11 DOWNTO 2);
			WHEN 519 => temp(5199 DOWNTO 5190) := ADC(11 DOWNTO 2);
			WHEN 520 => temp(5209 DOWNTO 5200) := ADC(11 DOWNTO 2);
			WHEN 521 => temp(5219 DOWNTO 5210) := ADC(11 DOWNTO 2);
			WHEN 522 => temp(5229 DOWNTO 5220) := ADC(11 DOWNTO 2);
			WHEN 523 => temp(5239 DOWNTO 5230) := ADC(11 DOWNTO 2);
			WHEN 524 => temp(5249 DOWNTO 5240) := ADC(11 DOWNTO 2);
			WHEN 525 => temp(5259 DOWNTO 5250) := ADC(11 DOWNTO 2);
			WHEN 526 => temp(5269 DOWNTO 5260) := ADC(11 DOWNTO 2);
			WHEN 527 => temp(5279 DOWNTO 5270) := ADC(11 DOWNTO 2);
			WHEN 528 => temp(5289 DOWNTO 5280) := ADC(11 DOWNTO 2);
			WHEN 529 => temp(5299 DOWNTO 5290) := ADC(11 DOWNTO 2);
			WHEN 530 => temp(5309 DOWNTO 5300) := ADC(11 DOWNTO 2);
			WHEN 531 => temp(5319 DOWNTO 5310) := ADC(11 DOWNTO 2);
			WHEN 532 => temp(5329 DOWNTO 5320) := ADC(11 DOWNTO 2);
			WHEN 533 => temp(5339 DOWNTO 5330) := ADC(11 DOWNTO 2);
			WHEN 534 => temp(5349 DOWNTO 5340) := ADC(11 DOWNTO 2);
			WHEN 535 => temp(5359 DOWNTO 5350) := ADC(11 DOWNTO 2);
			WHEN 536 => temp(5369 DOWNTO 5360) := ADC(11 DOWNTO 2);
			WHEN 537 => temp(5379 DOWNTO 5370) := ADC(11 DOWNTO 2);
			WHEN 538 => temp(5389 DOWNTO 5380) := ADC(11 DOWNTO 2);
			WHEN 539 => temp(5399 DOWNTO 5390) := ADC(11 DOWNTO 2);
			WHEN 540 => temp(5409 DOWNTO 5400) := ADC(11 DOWNTO 2);
			WHEN 541 => temp(5419 DOWNTO 5410) := ADC(11 DOWNTO 2);
			WHEN 542 => temp(5429 DOWNTO 5420) := ADC(11 DOWNTO 2);
			WHEN 543 => temp(5439 DOWNTO 5430) := ADC(11 DOWNTO 2);
			WHEN 544 => temp(5449 DOWNTO 5440) := ADC(11 DOWNTO 2);
			WHEN 545 => temp(5459 DOWNTO 5450) := ADC(11 DOWNTO 2);
			WHEN 546 => temp(5469 DOWNTO 5460) := ADC(11 DOWNTO 2);
			WHEN 547 => temp(5479 DOWNTO 5470) := ADC(11 DOWNTO 2);
			WHEN 548 => temp(5489 DOWNTO 5480) := ADC(11 DOWNTO 2);
			WHEN 549 => temp(5499 DOWNTO 5490) := ADC(11 DOWNTO 2);
			WHEN 550 => temp(5509 DOWNTO 5500) := ADC(11 DOWNTO 2);
			WHEN 551 => temp(5519 DOWNTO 5510) := ADC(11 DOWNTO 2);
			WHEN 552 => temp(5529 DOWNTO 5520) := ADC(11 DOWNTO 2);
			WHEN 553 => temp(5539 DOWNTO 5530) := ADC(11 DOWNTO 2);
			WHEN 554 => temp(5549 DOWNTO 5540) := ADC(11 DOWNTO 2);
			WHEN 555 => temp(5559 DOWNTO 5550) := ADC(11 DOWNTO 2);
			WHEN 556 => temp(5569 DOWNTO 5560) := ADC(11 DOWNTO 2);
			WHEN 557 => temp(5579 DOWNTO 5570) := ADC(11 DOWNTO 2);
			WHEN 558 => temp(5589 DOWNTO 5580) := ADC(11 DOWNTO 2);
			WHEN 559 => temp(5599 DOWNTO 5590) := ADC(11 DOWNTO 2);
			WHEN 560 => temp(5609 DOWNTO 5600) := ADC(11 DOWNTO 2);
			WHEN 561 => temp(5619 DOWNTO 5610) := ADC(11 DOWNTO 2);
			WHEN 562 => temp(5629 DOWNTO 5620) := ADC(11 DOWNTO 2);
			WHEN 563 => temp(5639 DOWNTO 5630) := ADC(11 DOWNTO 2);
			WHEN 564 => temp(5649 DOWNTO 5640) := ADC(11 DOWNTO 2);
			WHEN 565 => temp(5659 DOWNTO 5650) := ADC(11 DOWNTO 2);
			WHEN 566 => temp(5669 DOWNTO 5660) := ADC(11 DOWNTO 2);
			WHEN 567 => temp(5679 DOWNTO 5670) := ADC(11 DOWNTO 2);
			WHEN 568 => temp(5689 DOWNTO 5680) := ADC(11 DOWNTO 2);
			WHEN 569 => temp(5699 DOWNTO 5690) := ADC(11 DOWNTO 2);
			WHEN 570 => temp(5709 DOWNTO 5700) := ADC(11 DOWNTO 2);
			WHEN 571 => temp(5719 DOWNTO 5710) := ADC(11 DOWNTO 2);
			WHEN 572 => temp(5729 DOWNTO 5720) := ADC(11 DOWNTO 2);
			WHEN 573 => temp(5739 DOWNTO 5730) := ADC(11 DOWNTO 2);
			WHEN 574 => temp(5749 DOWNTO 5740) := ADC(11 DOWNTO 2);
			WHEN 575 => temp(5759 DOWNTO 5750) := ADC(11 DOWNTO 2);
			WHEN 576 => temp(5769 DOWNTO 5760) := ADC(11 DOWNTO 2);
			WHEN 577 => temp(5779 DOWNTO 5770) := ADC(11 DOWNTO 2);
			WHEN 578 => temp(5789 DOWNTO 5780) := ADC(11 DOWNTO 2);
			WHEN 579 => temp(5799 DOWNTO 5790) := ADC(11 DOWNTO 2);
			WHEN 580 => temp(5809 DOWNTO 5800) := ADC(11 DOWNTO 2);
			WHEN 581 => temp(5819 DOWNTO 5810) := ADC(11 DOWNTO 2);
			WHEN 582 => temp(5829 DOWNTO 5820) := ADC(11 DOWNTO 2);
			WHEN 583 => temp(5839 DOWNTO 5830) := ADC(11 DOWNTO 2);
			WHEN 584 => temp(5849 DOWNTO 5840) := ADC(11 DOWNTO 2);
			WHEN 585 => temp(5859 DOWNTO 5850) := ADC(11 DOWNTO 2);
			WHEN 586 => temp(5869 DOWNTO 5860) := ADC(11 DOWNTO 2);
			WHEN 587 => temp(5879 DOWNTO 5870) := ADC(11 DOWNTO 2);
			WHEN 588 => temp(5889 DOWNTO 5880) := ADC(11 DOWNTO 2);
			WHEN 589 => temp(5899 DOWNTO 5890) := ADC(11 DOWNTO 2);
			WHEN 590 => temp(5909 DOWNTO 5900) := ADC(11 DOWNTO 2);
			WHEN 591 => temp(5919 DOWNTO 5910) := ADC(11 DOWNTO 2);
			WHEN 592 => temp(5929 DOWNTO 5920) := ADC(11 DOWNTO 2);
			WHEN 593 => temp(5939 DOWNTO 5930) := ADC(11 DOWNTO 2);
			WHEN 594 => temp(5949 DOWNTO 5940) := ADC(11 DOWNTO 2);
			WHEN 595 => temp(5959 DOWNTO 5950) := ADC(11 DOWNTO 2);
			WHEN 596 => temp(5969 DOWNTO 5960) := ADC(11 DOWNTO 2);
			WHEN 597 => temp(5979 DOWNTO 5970) := ADC(11 DOWNTO 2);
			WHEN 598 => temp(5989 DOWNTO 5980) := ADC(11 DOWNTO 2);
			WHEN 599 => temp(5999 DOWNTO 5990) := ADC(11 DOWNTO 2);
			WHEN 600 => temp(6009 DOWNTO 6000) := ADC(11 DOWNTO 2);
			WHEN 601 => temp(6019 DOWNTO 6010) := ADC(11 DOWNTO 2);
			WHEN 602 => temp(6029 DOWNTO 6020) := ADC(11 DOWNTO 2);
			WHEN 603 => temp(6039 DOWNTO 6030) := ADC(11 DOWNTO 2);
			WHEN 604 => temp(6049 DOWNTO 6040) := ADC(11 DOWNTO 2);
			WHEN 605 => temp(6059 DOWNTO 6050) := ADC(11 DOWNTO 2);
			WHEN 606 => temp(6069 DOWNTO 6060) := ADC(11 DOWNTO 2);
			WHEN 607 => temp(6079 DOWNTO 6070) := ADC(11 DOWNTO 2);
			WHEN 608 => temp(6089 DOWNTO 6080) := ADC(11 DOWNTO 2);
			WHEN 609 => temp(6099 DOWNTO 6090) := ADC(11 DOWNTO 2);
			WHEN 610 => temp(6109 DOWNTO 6100) := ADC(11 DOWNTO 2);
			WHEN 611 => temp(6119 DOWNTO 6110) := ADC(11 DOWNTO 2);
			WHEN 612 => temp(6129 DOWNTO 6120) := ADC(11 DOWNTO 2);
			WHEN 613 => temp(6139 DOWNTO 6130) := ADC(11 DOWNTO 2);
			WHEN 614 => temp(6149 DOWNTO 6140) := ADC(11 DOWNTO 2);
			WHEN 615 => temp(6159 DOWNTO 6150) := ADC(11 DOWNTO 2);
			WHEN 616 => temp(6169 DOWNTO 6160) := ADC(11 DOWNTO 2);
			WHEN 617 => temp(6179 DOWNTO 6170) := ADC(11 DOWNTO 2);
			WHEN 618 => temp(6189 DOWNTO 6180) := ADC(11 DOWNTO 2);
			WHEN 619 => temp(6199 DOWNTO 6190) := ADC(11 DOWNTO 2);
			WHEN 620 => temp(6209 DOWNTO 6200) := ADC(11 DOWNTO 2);
			WHEN 621 => temp(6219 DOWNTO 6210) := ADC(11 DOWNTO 2);
			WHEN 622 => temp(6229 DOWNTO 6220) := ADC(11 DOWNTO 2);
			WHEN 623 => temp(6239 DOWNTO 6230) := ADC(11 DOWNTO 2);
			WHEN 624 => temp(6249 DOWNTO 6240) := ADC(11 DOWNTO 2);
			WHEN 625 => temp(6259 DOWNTO 6250) := ADC(11 DOWNTO 2);
			WHEN 626 => temp(6269 DOWNTO 6260) := ADC(11 DOWNTO 2);
			WHEN 627 => temp(6279 DOWNTO 6270) := ADC(11 DOWNTO 2);
			WHEN 628 => temp(6289 DOWNTO 6280) := ADC(11 DOWNTO 2);
			WHEN 629 => temp(6299 DOWNTO 6290) := ADC(11 DOWNTO 2);
			WHEN 630 => temp(6309 DOWNTO 6300) := ADC(11 DOWNTO 2);
			WHEN 631 => temp(6319 DOWNTO 6310) := ADC(11 DOWNTO 2);
			WHEN 632 => temp(6329 DOWNTO 6320) := ADC(11 DOWNTO 2);
			WHEN 633 => temp(6339 DOWNTO 6330) := ADC(11 DOWNTO 2);
			WHEN 634 => temp(6349 DOWNTO 6340) := ADC(11 DOWNTO 2);
			WHEN 635 => temp(6359 DOWNTO 6350) := ADC(11 DOWNTO 2);
			WHEN 636 => temp(6369 DOWNTO 6360) := ADC(11 DOWNTO 2);
			WHEN 637 => temp(6379 DOWNTO 6370) := ADC(11 DOWNTO 2);
			WHEN 638 => temp(6389 DOWNTO 6380) := ADC(11 DOWNTO 2);
			WHEN 639 => temp(6399 DOWNTO 6390) := ADC(11 DOWNTO 2);
			WHEN 640 => temp(6409 DOWNTO 6400) := ADC(11 DOWNTO 2);
			WHEN 641 => temp(6419 DOWNTO 6410) := ADC(11 DOWNTO 2);
			WHEN 642 => temp(6429 DOWNTO 6420) := ADC(11 DOWNTO 2);
			WHEN 643 => temp(6439 DOWNTO 6430) := ADC(11 DOWNTO 2);
			WHEN 644 => temp(6449 DOWNTO 6440) := ADC(11 DOWNTO 2);
			WHEN 645 => temp(6459 DOWNTO 6450) := ADC(11 DOWNTO 2);
			WHEN 646 => temp(6469 DOWNTO 6460) := ADC(11 DOWNTO 2);
			WHEN 647 => temp(6479 DOWNTO 6470) := ADC(11 DOWNTO 2);
			WHEN 648 => temp(6489 DOWNTO 6480) := ADC(11 DOWNTO 2);
			WHEN 649 => temp(6499 DOWNTO 6490) := ADC(11 DOWNTO 2);
			WHEN 650 => temp(6509 DOWNTO 6500) := ADC(11 DOWNTO 2);
			WHEN 651 => temp(6519 DOWNTO 6510) := ADC(11 DOWNTO 2);
			WHEN 652 => temp(6529 DOWNTO 6520) := ADC(11 DOWNTO 2);
			WHEN 653 => temp(6539 DOWNTO 6530) := ADC(11 DOWNTO 2);
			WHEN 654 => temp(6549 DOWNTO 6540) := ADC(11 DOWNTO 2);
			WHEN 655 => temp(6559 DOWNTO 6550) := ADC(11 DOWNTO 2);
			WHEN 656 => temp(6569 DOWNTO 6560) := ADC(11 DOWNTO 2);
			WHEN 657 => temp(6579 DOWNTO 6570) := ADC(11 DOWNTO 2);
			WHEN 658 => temp(6589 DOWNTO 6580) := ADC(11 DOWNTO 2);
			WHEN 659 => temp(6599 DOWNTO 6590) := ADC(11 DOWNTO 2);
			WHEN 660 => temp(6609 DOWNTO 6600) := ADC(11 DOWNTO 2);
			WHEN 661 => temp(6619 DOWNTO 6610) := ADC(11 DOWNTO 2);
			WHEN 662 => temp(6629 DOWNTO 6620) := ADC(11 DOWNTO 2);
			WHEN 663 => temp(6639 DOWNTO 6630) := ADC(11 DOWNTO 2);
			WHEN 664 => temp(6649 DOWNTO 6640) := ADC(11 DOWNTO 2);
			WHEN 665 => temp(6659 DOWNTO 6650) := ADC(11 DOWNTO 2);
			WHEN 666 => temp(6669 DOWNTO 6660) := ADC(11 DOWNTO 2);
			WHEN 667 => temp(6679 DOWNTO 6670) := ADC(11 DOWNTO 2);
			WHEN 668 => temp(6689 DOWNTO 6680) := ADC(11 DOWNTO 2);
			WHEN 669 => temp(6699 DOWNTO 6690) := ADC(11 DOWNTO 2);
			WHEN 670 => temp(6709 DOWNTO 6700) := ADC(11 DOWNTO 2);
			WHEN 671 => temp(6719 DOWNTO 6710) := ADC(11 DOWNTO 2);
			WHEN 672 => temp(6729 DOWNTO 6720) := ADC(11 DOWNTO 2);
			WHEN 673 => temp(6739 DOWNTO 6730) := ADC(11 DOWNTO 2);
			WHEN 674 => temp(6749 DOWNTO 6740) := ADC(11 DOWNTO 2);
			WHEN 675 => temp(6759 DOWNTO 6750) := ADC(11 DOWNTO 2);
			WHEN 676 => temp(6769 DOWNTO 6760) := ADC(11 DOWNTO 2);
			WHEN 677 => temp(6779 DOWNTO 6770) := ADC(11 DOWNTO 2);
			WHEN 678 => temp(6789 DOWNTO 6780) := ADC(11 DOWNTO 2);
			WHEN 679 => temp(6799 DOWNTO 6790) := ADC(11 DOWNTO 2);
			WHEN 680 => temp(6809 DOWNTO 6800) := ADC(11 DOWNTO 2);
			WHEN 681 => temp(6819 DOWNTO 6810) := ADC(11 DOWNTO 2);
			WHEN 682 => temp(6829 DOWNTO 6820) := ADC(11 DOWNTO 2);
			WHEN 683 => temp(6839 DOWNTO 6830) := ADC(11 DOWNTO 2);
			WHEN 684 => temp(6849 DOWNTO 6840) := ADC(11 DOWNTO 2);
			WHEN 685 => temp(6859 DOWNTO 6850) := ADC(11 DOWNTO 2);
			WHEN 686 => temp(6869 DOWNTO 6860) := ADC(11 DOWNTO 2);
			WHEN 687 => temp(6879 DOWNTO 6870) := ADC(11 DOWNTO 2);
			WHEN 688 => temp(6889 DOWNTO 6880) := ADC(11 DOWNTO 2);
			WHEN 689 => temp(6899 DOWNTO 6890) := ADC(11 DOWNTO 2);
			WHEN 690 => temp(6909 DOWNTO 6900) := ADC(11 DOWNTO 2);
			WHEN 691 => temp(6919 DOWNTO 6910) := ADC(11 DOWNTO 2);
			WHEN 692 => temp(6929 DOWNTO 6920) := ADC(11 DOWNTO 2);
			WHEN 693 => temp(6939 DOWNTO 6930) := ADC(11 DOWNTO 2);
			WHEN 694 => temp(6949 DOWNTO 6940) := ADC(11 DOWNTO 2);
			WHEN 695 => temp(6959 DOWNTO 6950) := ADC(11 DOWNTO 2);
			WHEN 696 => temp(6969 DOWNTO 6960) := ADC(11 DOWNTO 2);
			WHEN 697 => temp(6979 DOWNTO 6970) := ADC(11 DOWNTO 2);
			WHEN 698 => temp(6989 DOWNTO 6980) := ADC(11 DOWNTO 2);
			WHEN 699 => temp(6999 DOWNTO 6990) := ADC(11 DOWNTO 2);
			WHEN 700 => temp(7009 DOWNTO 7000) := ADC(11 DOWNTO 2);
			WHEN 701 => temp(7019 DOWNTO 7010) := ADC(11 DOWNTO 2);
			WHEN 702 => temp(7029 DOWNTO 7020) := ADC(11 DOWNTO 2);
			WHEN 703 => temp(7039 DOWNTO 7030) := ADC(11 DOWNTO 2);
			WHEN 704 => temp(7049 DOWNTO 7040) := ADC(11 DOWNTO 2);
			WHEN 705 => temp(7059 DOWNTO 7050) := ADC(11 DOWNTO 2);
			WHEN 706 => temp(7069 DOWNTO 7060) := ADC(11 DOWNTO 2);
			WHEN 707 => temp(7079 DOWNTO 7070) := ADC(11 DOWNTO 2);
			WHEN 708 => temp(7089 DOWNTO 7080) := ADC(11 DOWNTO 2);
			WHEN 709 => temp(7099 DOWNTO 7090) := ADC(11 DOWNTO 2);
			WHEN 710 => temp(7109 DOWNTO 7100) := ADC(11 DOWNTO 2);
			WHEN 711 => temp(7119 DOWNTO 7110) := ADC(11 DOWNTO 2);
			WHEN 712 => temp(7129 DOWNTO 7120) := ADC(11 DOWNTO 2);
			WHEN 713 => temp(7139 DOWNTO 7130) := ADC(11 DOWNTO 2);
			WHEN 714 => temp(7149 DOWNTO 7140) := ADC(11 DOWNTO 2);
			WHEN 715 => temp(7159 DOWNTO 7150) := ADC(11 DOWNTO 2);
			WHEN 716 => temp(7169 DOWNTO 7160) := ADC(11 DOWNTO 2);
			WHEN 717 => temp(7179 DOWNTO 7170) := ADC(11 DOWNTO 2);
			WHEN 718 => temp(7189 DOWNTO 7180) := ADC(11 DOWNTO 2);
			WHEN 719 => temp(7199 DOWNTO 7190) := ADC(11 DOWNTO 2);
			WHEN 720 => temp(7209 DOWNTO 7200) := ADC(11 DOWNTO 2);
			WHEN 721 => temp(7219 DOWNTO 7210) := ADC(11 DOWNTO 2);
			WHEN 722 => temp(7229 DOWNTO 7220) := ADC(11 DOWNTO 2);
			WHEN 723 => temp(7239 DOWNTO 7230) := ADC(11 DOWNTO 2);
			WHEN 724 => temp(7249 DOWNTO 7240) := ADC(11 DOWNTO 2);
			WHEN 725 => temp(7259 DOWNTO 7250) := ADC(11 DOWNTO 2);
			WHEN 726 => temp(7269 DOWNTO 7260) := ADC(11 DOWNTO 2);
			WHEN 727 => temp(7279 DOWNTO 7270) := ADC(11 DOWNTO 2);
			WHEN 728 => temp(7289 DOWNTO 7280) := ADC(11 DOWNTO 2);
			WHEN 729 => temp(7299 DOWNTO 7290) := ADC(11 DOWNTO 2);
			WHEN 730 => temp(7309 DOWNTO 7300) := ADC(11 DOWNTO 2);
			WHEN 731 => temp(7319 DOWNTO 7310) := ADC(11 DOWNTO 2);
			WHEN 732 => temp(7329 DOWNTO 7320) := ADC(11 DOWNTO 2);
			WHEN 733 => temp(7339 DOWNTO 7330) := ADC(11 DOWNTO 2);
			WHEN 734 => temp(7349 DOWNTO 7340) := ADC(11 DOWNTO 2);
			WHEN 735 => temp(7359 DOWNTO 7350) := ADC(11 DOWNTO 2);
			WHEN 736 => temp(7369 DOWNTO 7360) := ADC(11 DOWNTO 2);
			WHEN 737 => temp(7379 DOWNTO 7370) := ADC(11 DOWNTO 2);
			WHEN 738 => temp(7389 DOWNTO 7380) := ADC(11 DOWNTO 2);
			WHEN 739 => temp(7399 DOWNTO 7390) := ADC(11 DOWNTO 2);
			WHEN 740 => temp(7409 DOWNTO 7400) := ADC(11 DOWNTO 2);
			WHEN 741 => temp(7419 DOWNTO 7410) := ADC(11 DOWNTO 2);
			WHEN 742 => temp(7429 DOWNTO 7420) := ADC(11 DOWNTO 2);
			WHEN 743 => temp(7439 DOWNTO 7430) := ADC(11 DOWNTO 2);
			WHEN 744 => temp(7449 DOWNTO 7440) := ADC(11 DOWNTO 2);
			WHEN 745 => temp(7459 DOWNTO 7450) := ADC(11 DOWNTO 2);
			WHEN 746 => temp(7469 DOWNTO 7460) := ADC(11 DOWNTO 2);
			WHEN 747 => temp(7479 DOWNTO 7470) := ADC(11 DOWNTO 2);
			WHEN 748 => temp(7489 DOWNTO 7480) := ADC(11 DOWNTO 2);
			WHEN 749 => temp(7499 DOWNTO 7490) := ADC(11 DOWNTO 2);
			WHEN 750 => temp(7509 DOWNTO 7500) := ADC(11 DOWNTO 2);
			WHEN 751 => temp(7519 DOWNTO 7510) := ADC(11 DOWNTO 2);
			WHEN 752 => temp(7529 DOWNTO 7520) := ADC(11 DOWNTO 2);
			WHEN 753 => temp(7539 DOWNTO 7530) := ADC(11 DOWNTO 2);
			WHEN 754 => temp(7549 DOWNTO 7540) := ADC(11 DOWNTO 2);
			WHEN 755 => temp(7559 DOWNTO 7550) := ADC(11 DOWNTO 2);
			WHEN 756 => temp(7569 DOWNTO 7560) := ADC(11 DOWNTO 2);
			WHEN 757 => temp(7579 DOWNTO 7570) := ADC(11 DOWNTO 2);
			WHEN 758 => temp(7589 DOWNTO 7580) := ADC(11 DOWNTO 2);
			WHEN 759 => temp(7599 DOWNTO 7590) := ADC(11 DOWNTO 2);
			WHEN 760 => temp(7609 DOWNTO 7600) := ADC(11 DOWNTO 2);
			WHEN 761 => temp(7619 DOWNTO 7610) := ADC(11 DOWNTO 2);
			WHEN 762 => temp(7629 DOWNTO 7620) := ADC(11 DOWNTO 2);
			WHEN 763 => temp(7639 DOWNTO 7630) := ADC(11 DOWNTO 2);
			WHEN 764 => temp(7649 DOWNTO 7640) := ADC(11 DOWNTO 2);
			WHEN 765 => temp(7659 DOWNTO 7650) := ADC(11 DOWNTO 2);
			WHEN 766 => temp(7669 DOWNTO 7660) := ADC(11 DOWNTO 2);
			WHEN 767 => temp(7679 DOWNTO 7670) := ADC(11 DOWNTO 2);
			WHEN 768 => temp(7689 DOWNTO 7680) := ADC(11 DOWNTO 2);
			WHEN 769 => temp(7699 DOWNTO 7690) := ADC(11 DOWNTO 2);
			WHEN 770 => temp(7709 DOWNTO 7700) := ADC(11 DOWNTO 2);
			WHEN 771 => temp(7719 DOWNTO 7710) := ADC(11 DOWNTO 2);
			WHEN 772 => temp(7729 DOWNTO 7720) := ADC(11 DOWNTO 2);
			WHEN 773 => temp(7739 DOWNTO 7730) := ADC(11 DOWNTO 2);
			WHEN 774 => temp(7749 DOWNTO 7740) := ADC(11 DOWNTO 2);
			WHEN 775 => temp(7759 DOWNTO 7750) := ADC(11 DOWNTO 2);
			WHEN 776 => temp(7769 DOWNTO 7760) := ADC(11 DOWNTO 2);
			WHEN 777 => temp(7779 DOWNTO 7770) := ADC(11 DOWNTO 2);
			WHEN 778 => temp(7789 DOWNTO 7780) := ADC(11 DOWNTO 2);
			WHEN 779 => temp(7799 DOWNTO 7790) := ADC(11 DOWNTO 2);
			WHEN 780 => temp(7809 DOWNTO 7800) := ADC(11 DOWNTO 2);
			WHEN 781 => temp(7819 DOWNTO 7810) := ADC(11 DOWNTO 2);
			WHEN 782 => temp(7829 DOWNTO 7820) := ADC(11 DOWNTO 2);
			WHEN 783 => temp(7839 DOWNTO 7830) := ADC(11 DOWNTO 2);
			WHEN 784 => temp(7849 DOWNTO 7840) := ADC(11 DOWNTO 2);
			WHEN 785 => temp(7859 DOWNTO 7850) := ADC(11 DOWNTO 2);
			WHEN 786 => temp(7869 DOWNTO 7860) := ADC(11 DOWNTO 2);
			WHEN 787 => temp(7879 DOWNTO 7870) := ADC(11 DOWNTO 2);
			WHEN 788 => temp(7889 DOWNTO 7880) := ADC(11 DOWNTO 2);
			WHEN 789 => temp(7899 DOWNTO 7890) := ADC(11 DOWNTO 2);
			WHEN 790 => temp(7909 DOWNTO 7900) := ADC(11 DOWNTO 2);
			WHEN 791 => temp(7919 DOWNTO 7910) := ADC(11 DOWNTO 2);
			WHEN 792 => temp(7929 DOWNTO 7920) := ADC(11 DOWNTO 2);
			WHEN 793 => temp(7939 DOWNTO 7930) := ADC(11 DOWNTO 2);
			WHEN 794 => temp(7949 DOWNTO 7940) := ADC(11 DOWNTO 2);
			WHEN 795 => temp(7959 DOWNTO 7950) := ADC(11 DOWNTO 2);
			WHEN 796 => temp(7969 DOWNTO 7960) := ADC(11 DOWNTO 2);
			WHEN 797 => temp(7979 DOWNTO 7970) := ADC(11 DOWNTO 2);
			WHEN 798 => temp(7989 DOWNTO 7980) := ADC(11 DOWNTO 2);
			WHEN 799 => temp(7999 DOWNTO 7990) := ADC(11 DOWNTO 2);
			WHEN 800 => temp(8009 DOWNTO 8000) := ADC(11 DOWNTO 2);
			WHEN 801 => temp(8019 DOWNTO 8010) := ADC(11 DOWNTO 2);
			WHEN 802 => temp(8029 DOWNTO 8020) := ADC(11 DOWNTO 2);
			WHEN 803 => temp(8039 DOWNTO 8030) := ADC(11 DOWNTO 2);
			WHEN 804 => temp(8049 DOWNTO 8040) := ADC(11 DOWNTO 2);
			WHEN 805 => temp(8059 DOWNTO 8050) := ADC(11 DOWNTO 2);
			WHEN 806 => temp(8069 DOWNTO 8060) := ADC(11 DOWNTO 2);
			WHEN 807 => temp(8079 DOWNTO 8070) := ADC(11 DOWNTO 2);
			WHEN 808 => temp(8089 DOWNTO 8080) := ADC(11 DOWNTO 2);
			WHEN 809 => temp(8099 DOWNTO 8090) := ADC(11 DOWNTO 2);
			WHEN 810 => temp(8109 DOWNTO 8100) := ADC(11 DOWNTO 2);
			WHEN 811 => temp(8119 DOWNTO 8110) := ADC(11 DOWNTO 2);
			WHEN 812 => temp(8129 DOWNTO 8120) := ADC(11 DOWNTO 2);
			WHEN 813 => temp(8139 DOWNTO 8130) := ADC(11 DOWNTO 2);
			WHEN 814 => temp(8149 DOWNTO 8140) := ADC(11 DOWNTO 2);
			WHEN 815 => temp(8159 DOWNTO 8150) := ADC(11 DOWNTO 2);
			WHEN 816 => temp(8169 DOWNTO 8160) := ADC(11 DOWNTO 2);
			WHEN 817 => temp(8179 DOWNTO 8170) := ADC(11 DOWNTO 2);
			WHEN 818 => temp(8189 DOWNTO 8180) := ADC(11 DOWNTO 2);
			WHEN 819 => temp(8199 DOWNTO 8190) := ADC(11 DOWNTO 2);
			WHEN 820 => temp(8209 DOWNTO 8200) := ADC(11 DOWNTO 2);
			WHEN 821 => temp(8219 DOWNTO 8210) := ADC(11 DOWNTO 2);
			WHEN 822 => temp(8229 DOWNTO 8220) := ADC(11 DOWNTO 2);
			WHEN 823 => temp(8239 DOWNTO 8230) := ADC(11 DOWNTO 2);
			WHEN 824 => temp(8249 DOWNTO 8240) := ADC(11 DOWNTO 2);
			WHEN 825 => temp(8259 DOWNTO 8250) := ADC(11 DOWNTO 2);
			WHEN 826 => temp(8269 DOWNTO 8260) := ADC(11 DOWNTO 2);
			WHEN 827 => temp(8279 DOWNTO 8270) := ADC(11 DOWNTO 2);
			WHEN 828 => temp(8289 DOWNTO 8280) := ADC(11 DOWNTO 2);
			WHEN 829 => temp(8299 DOWNTO 8290) := ADC(11 DOWNTO 2);
			WHEN 830 => temp(8309 DOWNTO 8300) := ADC(11 DOWNTO 2);
			WHEN 831 => temp(8319 DOWNTO 8310) := ADC(11 DOWNTO 2);
			WHEN 832 => temp(8329 DOWNTO 8320) := ADC(11 DOWNTO 2);
			WHEN 833 => temp(8339 DOWNTO 8330) := ADC(11 DOWNTO 2);
			WHEN 834 => temp(8349 DOWNTO 8340) := ADC(11 DOWNTO 2);
			WHEN 835 => temp(8359 DOWNTO 8350) := ADC(11 DOWNTO 2);
			WHEN 836 => temp(8369 DOWNTO 8360) := ADC(11 DOWNTO 2);
			WHEN 837 => temp(8379 DOWNTO 8370) := ADC(11 DOWNTO 2);
			WHEN 838 => temp(8389 DOWNTO 8380) := ADC(11 DOWNTO 2);
			WHEN 839 => temp(8399 DOWNTO 8390) := ADC(11 DOWNTO 2);
			WHEN 840 => temp(8409 DOWNTO 8400) := ADC(11 DOWNTO 2);
			WHEN 841 => temp(8419 DOWNTO 8410) := ADC(11 DOWNTO 2);
			WHEN 842 => temp(8429 DOWNTO 8420) := ADC(11 DOWNTO 2);
			WHEN 843 => temp(8439 DOWNTO 8430) := ADC(11 DOWNTO 2);
			WHEN 844 => temp(8449 DOWNTO 8440) := ADC(11 DOWNTO 2);
			WHEN 845 => temp(8459 DOWNTO 8450) := ADC(11 DOWNTO 2);
			WHEN 846 => temp(8469 DOWNTO 8460) := ADC(11 DOWNTO 2);
			WHEN 847 => temp(8479 DOWNTO 8470) := ADC(11 DOWNTO 2);
			WHEN 848 => temp(8489 DOWNTO 8480) := ADC(11 DOWNTO 2);
			WHEN 849 => temp(8499 DOWNTO 8490) := ADC(11 DOWNTO 2);
			WHEN 850 => temp(8509 DOWNTO 8500) := ADC(11 DOWNTO 2);
			WHEN 851 => temp(8519 DOWNTO 8510) := ADC(11 DOWNTO 2);
			WHEN 852 => temp(8529 DOWNTO 8520) := ADC(11 DOWNTO 2);
			WHEN 853 => temp(8539 DOWNTO 8530) := ADC(11 DOWNTO 2);
			WHEN 854 => temp(8549 DOWNTO 8540) := ADC(11 DOWNTO 2);
			WHEN 855 => temp(8559 DOWNTO 8550) := ADC(11 DOWNTO 2);
			WHEN 856 => temp(8569 DOWNTO 8560) := ADC(11 DOWNTO 2);
			WHEN 857 => temp(8579 DOWNTO 8570) := ADC(11 DOWNTO 2);
			WHEN 858 => temp(8589 DOWNTO 8580) := ADC(11 DOWNTO 2);
			WHEN 859 => temp(8599 DOWNTO 8590) := ADC(11 DOWNTO 2);
			WHEN 860 => temp(8609 DOWNTO 8600) := ADC(11 DOWNTO 2);
			WHEN 861 => temp(8619 DOWNTO 8610) := ADC(11 DOWNTO 2);
			WHEN 862 => temp(8629 DOWNTO 8620) := ADC(11 DOWNTO 2);
			WHEN 863 => temp(8639 DOWNTO 8630) := ADC(11 DOWNTO 2);
			WHEN 864 => temp(8649 DOWNTO 8640) := ADC(11 DOWNTO 2);
			WHEN 865 => temp(8659 DOWNTO 8650) := ADC(11 DOWNTO 2);
			WHEN 866 => temp(8669 DOWNTO 8660) := ADC(11 DOWNTO 2);
			WHEN 867 => temp(8679 DOWNTO 8670) := ADC(11 DOWNTO 2);
			WHEN 868 => temp(8689 DOWNTO 8680) := ADC(11 DOWNTO 2);
			WHEN 869 => temp(8699 DOWNTO 8690) := ADC(11 DOWNTO 2);
			WHEN 870 => temp(8709 DOWNTO 8700) := ADC(11 DOWNTO 2);
			WHEN 871 => temp(8719 DOWNTO 8710) := ADC(11 DOWNTO 2);
			WHEN 872 => temp(8729 DOWNTO 8720) := ADC(11 DOWNTO 2);
			WHEN 873 => temp(8739 DOWNTO 8730) := ADC(11 DOWNTO 2);
			WHEN 874 => temp(8749 DOWNTO 8740) := ADC(11 DOWNTO 2);
			WHEN 875 => temp(8759 DOWNTO 8750) := ADC(11 DOWNTO 2);
			WHEN 876 => temp(8769 DOWNTO 8760) := ADC(11 DOWNTO 2);
			WHEN 877 => temp(8779 DOWNTO 8770) := ADC(11 DOWNTO 2);
			WHEN 878 => temp(8789 DOWNTO 8780) := ADC(11 DOWNTO 2);
			WHEN 879 => temp(8799 DOWNTO 8790) := ADC(11 DOWNTO 2);
			WHEN 880 => temp(8809 DOWNTO 8800) := ADC(11 DOWNTO 2);
			WHEN 881 => temp(8819 DOWNTO 8810) := ADC(11 DOWNTO 2);
			WHEN 882 => temp(8829 DOWNTO 8820) := ADC(11 DOWNTO 2);
			WHEN 883 => temp(8839 DOWNTO 8830) := ADC(11 DOWNTO 2);
			WHEN 884 => temp(8849 DOWNTO 8840) := ADC(11 DOWNTO 2);
			WHEN 885 => temp(8859 DOWNTO 8850) := ADC(11 DOWNTO 2);
			WHEN 886 => temp(8869 DOWNTO 8860) := ADC(11 DOWNTO 2);
			WHEN 887 => temp(8879 DOWNTO 8870) := ADC(11 DOWNTO 2);
			WHEN 888 => temp(8889 DOWNTO 8880) := ADC(11 DOWNTO 2);
			WHEN 889 => temp(8899 DOWNTO 8890) := ADC(11 DOWNTO 2);
			WHEN 890 => temp(8909 DOWNTO 8900) := ADC(11 DOWNTO 2);
			WHEN 891 => temp(8919 DOWNTO 8910) := ADC(11 DOWNTO 2);
			WHEN 892 => temp(8929 DOWNTO 8920) := ADC(11 DOWNTO 2);
			WHEN 893 => temp(8939 DOWNTO 8930) := ADC(11 DOWNTO 2);
			WHEN 894 => temp(8949 DOWNTO 8940) := ADC(11 DOWNTO 2);
			WHEN 895 => temp(8959 DOWNTO 8950) := ADC(11 DOWNTO 2);
			WHEN 896 => temp(8969 DOWNTO 8960) := ADC(11 DOWNTO 2);
			WHEN 897 => temp(8979 DOWNTO 8970) := ADC(11 DOWNTO 2);
			WHEN 898 => temp(8989 DOWNTO 8980) := ADC(11 DOWNTO 2);
			WHEN 899 => temp(8999 DOWNTO 8990) := ADC(11 DOWNTO 2);
			WHEN 900 => temp(9009 DOWNTO 9000) := ADC(11 DOWNTO 2);
			WHEN 901 => temp(9019 DOWNTO 9010) := ADC(11 DOWNTO 2);
			WHEN 902 => temp(9029 DOWNTO 9020) := ADC(11 DOWNTO 2);
			WHEN 903 => temp(9039 DOWNTO 9030) := ADC(11 DOWNTO 2);
			WHEN 904 => temp(9049 DOWNTO 9040) := ADC(11 DOWNTO 2);
			WHEN 905 => temp(9059 DOWNTO 9050) := ADC(11 DOWNTO 2);
			WHEN 906 => temp(9069 DOWNTO 9060) := ADC(11 DOWNTO 2);
			WHEN 907 => temp(9079 DOWNTO 9070) := ADC(11 DOWNTO 2);
			WHEN 908 => temp(9089 DOWNTO 9080) := ADC(11 DOWNTO 2);
			WHEN 909 => temp(9099 DOWNTO 9090) := ADC(11 DOWNTO 2);
			WHEN 910 => temp(9109 DOWNTO 9100) := ADC(11 DOWNTO 2);
			WHEN 911 => temp(9119 DOWNTO 9110) := ADC(11 DOWNTO 2);
			WHEN 912 => temp(9129 DOWNTO 9120) := ADC(11 DOWNTO 2);
			WHEN 913 => temp(9139 DOWNTO 9130) := ADC(11 DOWNTO 2);
			WHEN 914 => temp(9149 DOWNTO 9140) := ADC(11 DOWNTO 2);
			WHEN 915 => temp(9159 DOWNTO 9150) := ADC(11 DOWNTO 2);
			WHEN 916 => temp(9169 DOWNTO 9160) := ADC(11 DOWNTO 2);
			WHEN 917 => temp(9179 DOWNTO 9170) := ADC(11 DOWNTO 2);
			WHEN 918 => temp(9189 DOWNTO 9180) := ADC(11 DOWNTO 2);
			WHEN 919 => temp(9199 DOWNTO 9190) := ADC(11 DOWNTO 2);
			WHEN 920 => temp(9209 DOWNTO 9200) := ADC(11 DOWNTO 2);
			WHEN 921 => temp(9219 DOWNTO 9210) := ADC(11 DOWNTO 2);
			WHEN 922 => temp(9229 DOWNTO 9220) := ADC(11 DOWNTO 2);
			WHEN 923 => temp(9239 DOWNTO 9230) := ADC(11 DOWNTO 2);
			WHEN 924 => temp(9249 DOWNTO 9240) := ADC(11 DOWNTO 2);
			WHEN 925 => temp(9259 DOWNTO 9250) := ADC(11 DOWNTO 2);
			WHEN 926 => temp(9269 DOWNTO 9260) := ADC(11 DOWNTO 2);
			WHEN 927 => temp(9279 DOWNTO 9270) := ADC(11 DOWNTO 2);
			WHEN 928 => temp(9289 DOWNTO 9280) := ADC(11 DOWNTO 2);
			WHEN 929 => temp(9299 DOWNTO 9290) := ADC(11 DOWNTO 2);
			WHEN 930 => temp(9309 DOWNTO 9300) := ADC(11 DOWNTO 2);
			WHEN 931 => temp(9319 DOWNTO 9310) := ADC(11 DOWNTO 2);
			WHEN 932 => temp(9329 DOWNTO 9320) := ADC(11 DOWNTO 2);
			WHEN 933 => temp(9339 DOWNTO 9330) := ADC(11 DOWNTO 2);
			WHEN 934 => temp(9349 DOWNTO 9340) := ADC(11 DOWNTO 2);
			WHEN 935 => temp(9359 DOWNTO 9350) := ADC(11 DOWNTO 2);
			WHEN 936 => temp(9369 DOWNTO 9360) := ADC(11 DOWNTO 2);
			WHEN 937 => temp(9379 DOWNTO 9370) := ADC(11 DOWNTO 2);
			WHEN 938 => temp(9389 DOWNTO 9380) := ADC(11 DOWNTO 2);
			WHEN 939 => temp(9399 DOWNTO 9390) := ADC(11 DOWNTO 2);
			WHEN 940 => temp(9409 DOWNTO 9400) := ADC(11 DOWNTO 2);
			WHEN 941 => temp(9419 DOWNTO 9410) := ADC(11 DOWNTO 2);
			WHEN 942 => temp(9429 DOWNTO 9420) := ADC(11 DOWNTO 2);
			WHEN 943 => temp(9439 DOWNTO 9430) := ADC(11 DOWNTO 2);
			WHEN 944 => temp(9449 DOWNTO 9440) := ADC(11 DOWNTO 2);
			WHEN 945 => temp(9459 DOWNTO 9450) := ADC(11 DOWNTO 2);
			WHEN 946 => temp(9469 DOWNTO 9460) := ADC(11 DOWNTO 2);
			WHEN 947 => temp(9479 DOWNTO 9470) := ADC(11 DOWNTO 2);
			WHEN 948 => temp(9489 DOWNTO 9480) := ADC(11 DOWNTO 2);
			WHEN 949 => temp(9499 DOWNTO 9490) := ADC(11 DOWNTO 2);
			WHEN 950 => temp(9509 DOWNTO 9500) := ADC(11 DOWNTO 2);
			WHEN 951 => temp(9519 DOWNTO 9510) := ADC(11 DOWNTO 2);
			WHEN 952 => temp(9529 DOWNTO 9520) := ADC(11 DOWNTO 2);
			WHEN 953 => temp(9539 DOWNTO 9530) := ADC(11 DOWNTO 2);
			WHEN 954 => temp(9549 DOWNTO 9540) := ADC(11 DOWNTO 2);
			WHEN 955 => temp(9559 DOWNTO 9550) := ADC(11 DOWNTO 2);
			WHEN 956 => temp(9569 DOWNTO 9560) := ADC(11 DOWNTO 2);
			WHEN 957 => temp(9579 DOWNTO 9570) := ADC(11 DOWNTO 2);
			WHEN 958 => temp(9589 DOWNTO 9580) := ADC(11 DOWNTO 2);
			WHEN 959 => temp(9599 DOWNTO 9590) := ADC(11 DOWNTO 2);
			WHEN 960 => temp(9609 DOWNTO 9600) := ADC(11 DOWNTO 2);
			WHEN 961 => temp(9619 DOWNTO 9610) := ADC(11 DOWNTO 2);
			WHEN 962 => temp(9629 DOWNTO 9620) := ADC(11 DOWNTO 2);
			WHEN 963 => temp(9639 DOWNTO 9630) := ADC(11 DOWNTO 2);
			WHEN 964 => temp(9649 DOWNTO 9640) := ADC(11 DOWNTO 2);
			WHEN 965 => temp(9659 DOWNTO 9650) := ADC(11 DOWNTO 2);
			WHEN 966 => temp(9669 DOWNTO 9660) := ADC(11 DOWNTO 2);
			WHEN 967 => temp(9679 DOWNTO 9670) := ADC(11 DOWNTO 2);
			WHEN 968 => temp(9689 DOWNTO 9680) := ADC(11 DOWNTO 2);
			WHEN 969 => temp(9699 DOWNTO 9690) := ADC(11 DOWNTO 2);
			WHEN 970 => temp(9709 DOWNTO 9700) := ADC(11 DOWNTO 2);
			WHEN 971 => temp(9719 DOWNTO 9710) := ADC(11 DOWNTO 2);
			WHEN 972 => temp(9729 DOWNTO 9720) := ADC(11 DOWNTO 2);
			WHEN 973 => temp(9739 DOWNTO 9730) := ADC(11 DOWNTO 2);
			WHEN 974 => temp(9749 DOWNTO 9740) := ADC(11 DOWNTO 2);
			WHEN 975 => temp(9759 DOWNTO 9750) := ADC(11 DOWNTO 2);
			WHEN 976 => temp(9769 DOWNTO 9760) := ADC(11 DOWNTO 2);
			WHEN 977 => temp(9779 DOWNTO 9770) := ADC(11 DOWNTO 2);
			WHEN 978 => temp(9789 DOWNTO 9780) := ADC(11 DOWNTO 2);
			WHEN 979 => temp(9799 DOWNTO 9790) := ADC(11 DOWNTO 2);
			WHEN 980 => temp(9809 DOWNTO 9800) := ADC(11 DOWNTO 2);
			WHEN 981 => temp(9819 DOWNTO 9810) := ADC(11 DOWNTO 2);
			WHEN 982 => temp(9829 DOWNTO 9820) := ADC(11 DOWNTO 2);
			WHEN 983 => temp(9839 DOWNTO 9830) := ADC(11 DOWNTO 2);
			WHEN 984 => temp(9849 DOWNTO 9840) := ADC(11 DOWNTO 2);
			WHEN 985 => temp(9859 DOWNTO 9850) := ADC(11 DOWNTO 2);
			WHEN 986 => temp(9869 DOWNTO 9860) := ADC(11 DOWNTO 2);
			WHEN 987 => temp(9879 DOWNTO 9870) := ADC(11 DOWNTO 2);
			WHEN 988 => temp(9889 DOWNTO 9880) := ADC(11 DOWNTO 2);
			WHEN 989 => temp(9899 DOWNTO 9890) := ADC(11 DOWNTO 2);
			WHEN 990 => temp(9909 DOWNTO 9900) := ADC(11 DOWNTO 2);
			WHEN 991 => temp(9919 DOWNTO 9910) := ADC(11 DOWNTO 2);
			WHEN 992 => temp(9929 DOWNTO 9920) := ADC(11 DOWNTO 2);
			WHEN 993 => temp(9939 DOWNTO 9930) := ADC(11 DOWNTO 2);
			WHEN 994 => temp(9949 DOWNTO 9940) := ADC(11 DOWNTO 2);
			WHEN 995 => temp(9959 DOWNTO 9950) := ADC(11 DOWNTO 2);
			WHEN 996 => temp(9969 DOWNTO 9960) := ADC(11 DOWNTO 2);
			WHEN 997 => temp(9979 DOWNTO 9970) := ADC(11 DOWNTO 2);
			WHEN 998 => temp(9989 DOWNTO 9980) := ADC(11 DOWNTO 2);
			WHEN 999 => temp(9999 DOWNTO 9990) := ADC(11 DOWNTO 2);
			WHEN 1000 => temp(10009 DOWNTO 10000) := ADC(11 DOWNTO 2);
			WHEN 1001 => temp(10019 DOWNTO 10010) := ADC(11 DOWNTO 2);
			WHEN 1002 => temp(10029 DOWNTO 10020) := ADC(11 DOWNTO 2);
			WHEN 1003 => temp(10039 DOWNTO 10030) := ADC(11 DOWNTO 2);
			WHEN 1004 => temp(10049 DOWNTO 10040) := ADC(11 DOWNTO 2);
			WHEN 1005 => temp(10059 DOWNTO 10050) := ADC(11 DOWNTO 2);
			WHEN 1006 => temp(10069 DOWNTO 10060) := ADC(11 DOWNTO 2);
			WHEN 1007 => temp(10079 DOWNTO 10070) := ADC(11 DOWNTO 2);
			WHEN 1008 => temp(10089 DOWNTO 10080) := ADC(11 DOWNTO 2);
			WHEN 1009 => temp(10099 DOWNTO 10090) := ADC(11 DOWNTO 2);
			WHEN 1010 => temp(10109 DOWNTO 10100) := ADC(11 DOWNTO 2);
			WHEN 1011 => temp(10119 DOWNTO 10110) := ADC(11 DOWNTO 2);
			WHEN 1012 => temp(10129 DOWNTO 10120) := ADC(11 DOWNTO 2);
			WHEN 1013 => temp(10139 DOWNTO 10130) := ADC(11 DOWNTO 2);
			WHEN 1014 => temp(10149 DOWNTO 10140) := ADC(11 DOWNTO 2);
			WHEN 1015 => temp(10159 DOWNTO 10150) := ADC(11 DOWNTO 2);
			WHEN 1016 => temp(10169 DOWNTO 10160) := ADC(11 DOWNTO 2);
			WHEN 1017 => temp(10179 DOWNTO 10170) := ADC(11 DOWNTO 2);
			WHEN 1018 => temp(10189 DOWNTO 10180) := ADC(11 DOWNTO 2);
			WHEN 1019 => temp(10199 DOWNTO 10190) := ADC(11 DOWNTO 2);
			WHEN 1020 => temp(10209 DOWNTO 10200) := ADC(11 DOWNTO 2);
			WHEN 1021 => temp(10219 DOWNTO 10210) := ADC(11 DOWNTO 2);
			WHEN 1022 => temp(10229 DOWNTO 10220) := ADC(11 DOWNTO 2);
			WHEN 1023 => temp(10239 DOWNTO 10230) := ADC(11 DOWNTO 2);
			WHEN 1024 => temp(10249 DOWNTO 10240) := ADC(11 DOWNTO 2);
			WHEN 1025 => temp(10259 DOWNTO 10250) := ADC(11 DOWNTO 2);
			WHEN 1026 => temp(10269 DOWNTO 10260) := ADC(11 DOWNTO 2);
			WHEN 1027 => temp(10279 DOWNTO 10270) := ADC(11 DOWNTO 2);
			WHEN 1028 => temp(10289 DOWNTO 10280) := ADC(11 DOWNTO 2);
			WHEN 1029 => temp(10299 DOWNTO 10290) := ADC(11 DOWNTO 2);
			WHEN 1030 => temp(10309 DOWNTO 10300) := ADC(11 DOWNTO 2);
			WHEN 1031 => temp(10319 DOWNTO 10310) := ADC(11 DOWNTO 2);
			WHEN 1032 => temp(10329 DOWNTO 10320) := ADC(11 DOWNTO 2);
			WHEN 1033 => temp(10339 DOWNTO 10330) := ADC(11 DOWNTO 2);
			WHEN 1034 => temp(10349 DOWNTO 10340) := ADC(11 DOWNTO 2);
			WHEN 1035 => temp(10359 DOWNTO 10350) := ADC(11 DOWNTO 2);
			WHEN 1036 => temp(10369 DOWNTO 10360) := ADC(11 DOWNTO 2);
			WHEN 1037 => temp(10379 DOWNTO 10370) := ADC(11 DOWNTO 2);
			WHEN 1038 => temp(10389 DOWNTO 10380) := ADC(11 DOWNTO 2);
			WHEN 1039 => temp(10399 DOWNTO 10390) := ADC(11 DOWNTO 2);
			WHEN 1040 => temp(10409 DOWNTO 10400) := ADC(11 DOWNTO 2);
			WHEN 1041 => temp(10419 DOWNTO 10410) := ADC(11 DOWNTO 2);
			WHEN 1042 => temp(10429 DOWNTO 10420) := ADC(11 DOWNTO 2);
			WHEN 1043 => temp(10439 DOWNTO 10430) := ADC(11 DOWNTO 2);
			WHEN 1044 => temp(10449 DOWNTO 10440) := ADC(11 DOWNTO 2);
			WHEN 1045 => temp(10459 DOWNTO 10450) := ADC(11 DOWNTO 2);
			WHEN 1046 => temp(10469 DOWNTO 10460) := ADC(11 DOWNTO 2);
			WHEN 1047 => temp(10479 DOWNTO 10470) := ADC(11 DOWNTO 2);
			WHEN 1048 => temp(10489 DOWNTO 10480) := ADC(11 DOWNTO 2);
			WHEN 1049 => temp(10499 DOWNTO 10490) := ADC(11 DOWNTO 2);
			WHEN 1050 => temp(10509 DOWNTO 10500) := ADC(11 DOWNTO 2);
			WHEN 1051 => temp(10519 DOWNTO 10510) := ADC(11 DOWNTO 2);
			WHEN 1052 => temp(10529 DOWNTO 10520) := ADC(11 DOWNTO 2);
			WHEN 1053 => temp(10539 DOWNTO 10530) := ADC(11 DOWNTO 2);
			WHEN 1054 => temp(10549 DOWNTO 10540) := ADC(11 DOWNTO 2);
			WHEN 1055 => temp(10559 DOWNTO 10550) := ADC(11 DOWNTO 2);
			WHEN 1056 => temp(10569 DOWNTO 10560) := ADC(11 DOWNTO 2);
			WHEN 1057 => temp(10579 DOWNTO 10570) := ADC(11 DOWNTO 2);
			WHEN 1058 => temp(10589 DOWNTO 10580) := ADC(11 DOWNTO 2);
			WHEN 1059 => temp(10599 DOWNTO 10590) := ADC(11 DOWNTO 2);
			WHEN 1060 => temp(10609 DOWNTO 10600) := ADC(11 DOWNTO 2);
			WHEN 1061 => temp(10619 DOWNTO 10610) := ADC(11 DOWNTO 2);
			WHEN 1062 => temp(10629 DOWNTO 10620) := ADC(11 DOWNTO 2);
			WHEN 1063 => temp(10639 DOWNTO 10630) := ADC(11 DOWNTO 2);
			WHEN 1064 => temp(10649 DOWNTO 10640) := ADC(11 DOWNTO 2);
			WHEN 1065 => temp(10659 DOWNTO 10650) := ADC(11 DOWNTO 2);
			WHEN 1066 => temp(10669 DOWNTO 10660) := ADC(11 DOWNTO 2);
			WHEN 1067 => temp(10679 DOWNTO 10670) := ADC(11 DOWNTO 2);
			WHEN 1068 => temp(10689 DOWNTO 10680) := ADC(11 DOWNTO 2);
			WHEN 1069 => temp(10699 DOWNTO 10690) := ADC(11 DOWNTO 2);
			WHEN 1070 => temp(10709 DOWNTO 10700) := ADC(11 DOWNTO 2);
			WHEN 1071 => temp(10719 DOWNTO 10710) := ADC(11 DOWNTO 2);
			WHEN 1072 => temp(10729 DOWNTO 10720) := ADC(11 DOWNTO 2);
			WHEN 1073 => temp(10739 DOWNTO 10730) := ADC(11 DOWNTO 2);
			WHEN 1074 => temp(10749 DOWNTO 10740) := ADC(11 DOWNTO 2);
			WHEN 1075 => temp(10759 DOWNTO 10750) := ADC(11 DOWNTO 2);
			WHEN 1076 => temp(10769 DOWNTO 10760) := ADC(11 DOWNTO 2);
			WHEN 1077 => temp(10779 DOWNTO 10770) := ADC(11 DOWNTO 2);
			WHEN 1078 => temp(10789 DOWNTO 10780) := ADC(11 DOWNTO 2);
			WHEN 1079 => temp(10799 DOWNTO 10790) := ADC(11 DOWNTO 2);
			WHEN 1080 => temp(10809 DOWNTO 10800) := ADC(11 DOWNTO 2);
			WHEN 1081 => temp(10819 DOWNTO 10810) := ADC(11 DOWNTO 2);
			WHEN 1082 => temp(10829 DOWNTO 10820) := ADC(11 DOWNTO 2);
			WHEN 1083 => temp(10839 DOWNTO 10830) := ADC(11 DOWNTO 2);
			WHEN 1084 => temp(10849 DOWNTO 10840) := ADC(11 DOWNTO 2);
			WHEN 1085 => temp(10859 DOWNTO 10850) := ADC(11 DOWNTO 2);
			WHEN 1086 => temp(10869 DOWNTO 10860) := ADC(11 DOWNTO 2);
			WHEN 1087 => temp(10879 DOWNTO 10870) := ADC(11 DOWNTO 2);
			WHEN 1088 => temp(10889 DOWNTO 10880) := ADC(11 DOWNTO 2);
			WHEN 1089 => temp(10899 DOWNTO 10890) := ADC(11 DOWNTO 2);
			WHEN 1090 => temp(10909 DOWNTO 10900) := ADC(11 DOWNTO 2);
			WHEN 1091 => temp(10919 DOWNTO 10910) := ADC(11 DOWNTO 2);
			WHEN 1092 => temp(10929 DOWNTO 10920) := ADC(11 DOWNTO 2);
			WHEN 1093 => temp(10939 DOWNTO 10930) := ADC(11 DOWNTO 2);
			WHEN 1094 => temp(10949 DOWNTO 10940) := ADC(11 DOWNTO 2);
			WHEN 1095 => temp(10959 DOWNTO 10950) := ADC(11 DOWNTO 2);
			WHEN 1096 => temp(10969 DOWNTO 10960) := ADC(11 DOWNTO 2);
			WHEN 1097 => temp(10979 DOWNTO 10970) := ADC(11 DOWNTO 2);
			WHEN 1098 => temp(10989 DOWNTO 10980) := ADC(11 DOWNTO 2);
			WHEN 1099 => temp(10999 DOWNTO 10990) := ADC(11 DOWNTO 2);
			WHEN 1100 => temp(11009 DOWNTO 11000) := ADC(11 DOWNTO 2);
			WHEN 1101 => temp(11019 DOWNTO 11010) := ADC(11 DOWNTO 2);
			WHEN 1102 => temp(11029 DOWNTO 11020) := ADC(11 DOWNTO 2);
			WHEN 1103 => temp(11039 DOWNTO 11030) := ADC(11 DOWNTO 2);
			WHEN 1104 => temp(11049 DOWNTO 11040) := ADC(11 DOWNTO 2);
			WHEN 1105 => temp(11059 DOWNTO 11050) := ADC(11 DOWNTO 2);
			WHEN 1106 => temp(11069 DOWNTO 11060) := ADC(11 DOWNTO 2);
			WHEN 1107 => temp(11079 DOWNTO 11070) := ADC(11 DOWNTO 2);
			WHEN 1108 => temp(11089 DOWNTO 11080) := ADC(11 DOWNTO 2);
			WHEN 1109 => temp(11099 DOWNTO 11090) := ADC(11 DOWNTO 2);
			WHEN 1110 => temp(11109 DOWNTO 11100) := ADC(11 DOWNTO 2);
			WHEN 1111 => temp(11119 DOWNTO 11110) := ADC(11 DOWNTO 2);
			WHEN 1112 => temp(11129 DOWNTO 11120) := ADC(11 DOWNTO 2);
			WHEN 1113 => temp(11139 DOWNTO 11130) := ADC(11 DOWNTO 2);
			WHEN 1114 => temp(11149 DOWNTO 11140) := ADC(11 DOWNTO 2);
			WHEN 1115 => temp(11159 DOWNTO 11150) := ADC(11 DOWNTO 2);
			WHEN 1116 => temp(11169 DOWNTO 11160) := ADC(11 DOWNTO 2);
			WHEN 1117 => temp(11179 DOWNTO 11170) := ADC(11 DOWNTO 2);
			WHEN 1118 => temp(11189 DOWNTO 11180) := ADC(11 DOWNTO 2);
			WHEN 1119 => temp(11199 DOWNTO 11190) := ADC(11 DOWNTO 2);
			WHEN 1120 => temp(11209 DOWNTO 11200) := ADC(11 DOWNTO 2);
			WHEN 1121 => temp(11219 DOWNTO 11210) := ADC(11 DOWNTO 2);
			WHEN 1122 => temp(11229 DOWNTO 11220) := ADC(11 DOWNTO 2);
			WHEN 1123 => temp(11239 DOWNTO 11230) := ADC(11 DOWNTO 2);
			WHEN 1124 => temp(11249 DOWNTO 11240) := ADC(11 DOWNTO 2);
			WHEN 1125 => temp(11259 DOWNTO 11250) := ADC(11 DOWNTO 2);
			WHEN 1126 => temp(11269 DOWNTO 11260) := ADC(11 DOWNTO 2);
			WHEN 1127 => temp(11279 DOWNTO 11270) := ADC(11 DOWNTO 2);
			WHEN 1128 => temp(11289 DOWNTO 11280) := ADC(11 DOWNTO 2);
			WHEN 1129 => temp(11299 DOWNTO 11290) := ADC(11 DOWNTO 2);
			WHEN 1130 => temp(11309 DOWNTO 11300) := ADC(11 DOWNTO 2);
			WHEN 1131 => temp(11319 DOWNTO 11310) := ADC(11 DOWNTO 2);
			WHEN 1132 => temp(11329 DOWNTO 11320) := ADC(11 DOWNTO 2);
			WHEN 1133 => temp(11339 DOWNTO 11330) := ADC(11 DOWNTO 2);
			WHEN 1134 => temp(11349 DOWNTO 11340) := ADC(11 DOWNTO 2);
			WHEN 1135 => temp(11359 DOWNTO 11350) := ADC(11 DOWNTO 2);
			WHEN 1136 => temp(11369 DOWNTO 11360) := ADC(11 DOWNTO 2);
			WHEN 1137 => temp(11379 DOWNTO 11370) := ADC(11 DOWNTO 2);
			WHEN 1138 => temp(11389 DOWNTO 11380) := ADC(11 DOWNTO 2);
			WHEN 1139 => temp(11399 DOWNTO 11390) := ADC(11 DOWNTO 2);
			WHEN 1140 => temp(11409 DOWNTO 11400) := ADC(11 DOWNTO 2);
			WHEN 1141 => temp(11419 DOWNTO 11410) := ADC(11 DOWNTO 2);
			WHEN 1142 => temp(11429 DOWNTO 11420) := ADC(11 DOWNTO 2);
			WHEN 1143 => temp(11439 DOWNTO 11430) := ADC(11 DOWNTO 2);
			WHEN 1144 => temp(11449 DOWNTO 11440) := ADC(11 DOWNTO 2);
			WHEN 1145 => temp(11459 DOWNTO 11450) := ADC(11 DOWNTO 2);
			WHEN 1146 => temp(11469 DOWNTO 11460) := ADC(11 DOWNTO 2);
			WHEN 1147 => temp(11479 DOWNTO 11470) := ADC(11 DOWNTO 2);
			WHEN 1148 => temp(11489 DOWNTO 11480) := ADC(11 DOWNTO 2);
			WHEN 1149 => temp(11499 DOWNTO 11490) := ADC(11 DOWNTO 2);
			WHEN 1150 => temp(11509 DOWNTO 11500) := ADC(11 DOWNTO 2);
			WHEN 1151 => temp(11519 DOWNTO 11510) := ADC(11 DOWNTO 2);
			WHEN 1152 => temp(11529 DOWNTO 11520) := ADC(11 DOWNTO 2);
			WHEN 1153 => temp(11539 DOWNTO 11530) := ADC(11 DOWNTO 2);
			WHEN 1154 => temp(11549 DOWNTO 11540) := ADC(11 DOWNTO 2);
			WHEN 1155 => temp(11559 DOWNTO 11550) := ADC(11 DOWNTO 2);
			WHEN 1156 => temp(11569 DOWNTO 11560) := ADC(11 DOWNTO 2);
			WHEN 1157 => temp(11579 DOWNTO 11570) := ADC(11 DOWNTO 2);
			WHEN 1158 => temp(11589 DOWNTO 11580) := ADC(11 DOWNTO 2);
			WHEN 1159 => temp(11599 DOWNTO 11590) := ADC(11 DOWNTO 2);
			WHEN 1160 => temp(11609 DOWNTO 11600) := ADC(11 DOWNTO 2);
			WHEN 1161 => temp(11619 DOWNTO 11610) := ADC(11 DOWNTO 2);
			WHEN 1162 => temp(11629 DOWNTO 11620) := ADC(11 DOWNTO 2);
			WHEN 1163 => temp(11639 DOWNTO 11630) := ADC(11 DOWNTO 2);
			WHEN 1164 => temp(11649 DOWNTO 11640) := ADC(11 DOWNTO 2);
			WHEN 1165 => temp(11659 DOWNTO 11650) := ADC(11 DOWNTO 2);
			WHEN 1166 => temp(11669 DOWNTO 11660) := ADC(11 DOWNTO 2);
			WHEN 1167 => temp(11679 DOWNTO 11670) := ADC(11 DOWNTO 2);
			WHEN 1168 => temp(11689 DOWNTO 11680) := ADC(11 DOWNTO 2);
			WHEN 1169 => temp(11699 DOWNTO 11690) := ADC(11 DOWNTO 2);
			WHEN 1170 => temp(11709 DOWNTO 11700) := ADC(11 DOWNTO 2);
			WHEN 1171 => temp(11719 DOWNTO 11710) := ADC(11 DOWNTO 2);
			WHEN 1172 => temp(11729 DOWNTO 11720) := ADC(11 DOWNTO 2);
			WHEN 1173 => temp(11739 DOWNTO 11730) := ADC(11 DOWNTO 2);
			WHEN 1174 => temp(11749 DOWNTO 11740) := ADC(11 DOWNTO 2);
			WHEN 1175 => temp(11759 DOWNTO 11750) := ADC(11 DOWNTO 2);
			WHEN 1176 => temp(11769 DOWNTO 11760) := ADC(11 DOWNTO 2);
			WHEN 1177 => temp(11779 DOWNTO 11770) := ADC(11 DOWNTO 2);
			WHEN 1178 => temp(11789 DOWNTO 11780) := ADC(11 DOWNTO 2);
			WHEN 1179 => temp(11799 DOWNTO 11790) := ADC(11 DOWNTO 2);
			WHEN 1180 => temp(11809 DOWNTO 11800) := ADC(11 DOWNTO 2);
			WHEN 1181 => temp(11819 DOWNTO 11810) := ADC(11 DOWNTO 2);
			WHEN 1182 => temp(11829 DOWNTO 11820) := ADC(11 DOWNTO 2);
			WHEN 1183 => temp(11839 DOWNTO 11830) := ADC(11 DOWNTO 2);
			WHEN 1184 => temp(11849 DOWNTO 11840) := ADC(11 DOWNTO 2);
			WHEN 1185 => temp(11859 DOWNTO 11850) := ADC(11 DOWNTO 2);
			WHEN 1186 => temp(11869 DOWNTO 11860) := ADC(11 DOWNTO 2);
			WHEN 1187 => temp(11879 DOWNTO 11870) := ADC(11 DOWNTO 2);
			WHEN 1188 => temp(11889 DOWNTO 11880) := ADC(11 DOWNTO 2);
			WHEN 1189 => temp(11899 DOWNTO 11890) := ADC(11 DOWNTO 2);
			WHEN 1190 => temp(11909 DOWNTO 11900) := ADC(11 DOWNTO 2);
			WHEN 1191 => temp(11919 DOWNTO 11910) := ADC(11 DOWNTO 2);
			WHEN 1192 => temp(11929 DOWNTO 11920) := ADC(11 DOWNTO 2);
			WHEN 1193 => temp(11939 DOWNTO 11930) := ADC(11 DOWNTO 2);
			WHEN 1194 => temp(11949 DOWNTO 11940) := ADC(11 DOWNTO 2);
			WHEN 1195 => temp(11959 DOWNTO 11950) := ADC(11 DOWNTO 2);
			WHEN 1196 => temp(11969 DOWNTO 11960) := ADC(11 DOWNTO 2);
			WHEN 1197 => temp(11979 DOWNTO 11970) := ADC(11 DOWNTO 2);
			WHEN 1198 => temp(11989 DOWNTO 11980) := ADC(11 DOWNTO 2);
			WHEN 1199 => temp(11999 DOWNTO 11990) := ADC(11 DOWNTO 2);
			WHEN 1200 => temp(12009 DOWNTO 12000) := ADC(11 DOWNTO 2);
			WHEN 1201 => temp(12019 DOWNTO 12010) := ADC(11 DOWNTO 2);
			WHEN 1202 => temp(12029 DOWNTO 12020) := ADC(11 DOWNTO 2);
			WHEN 1203 => temp(12039 DOWNTO 12030) := ADC(11 DOWNTO 2);
			WHEN 1204 => temp(12049 DOWNTO 12040) := ADC(11 DOWNTO 2);
			WHEN 1205 => temp(12059 DOWNTO 12050) := ADC(11 DOWNTO 2);
			WHEN 1206 => temp(12069 DOWNTO 12060) := ADC(11 DOWNTO 2);
			WHEN 1207 => temp(12079 DOWNTO 12070) := ADC(11 DOWNTO 2);
			WHEN 1208 => temp(12089 DOWNTO 12080) := ADC(11 DOWNTO 2);
			WHEN 1209 => temp(12099 DOWNTO 12090) := ADC(11 DOWNTO 2);
			WHEN 1210 => temp(12109 DOWNTO 12100) := ADC(11 DOWNTO 2);
			WHEN 1211 => temp(12119 DOWNTO 12110) := ADC(11 DOWNTO 2);
			WHEN 1212 => temp(12129 DOWNTO 12120) := ADC(11 DOWNTO 2);
			WHEN 1213 => temp(12139 DOWNTO 12130) := ADC(11 DOWNTO 2);
			WHEN 1214 => temp(12149 DOWNTO 12140) := ADC(11 DOWNTO 2);
			WHEN 1215 => temp(12159 DOWNTO 12150) := ADC(11 DOWNTO 2);
			WHEN 1216 => temp(12169 DOWNTO 12160) := ADC(11 DOWNTO 2);
			WHEN 1217 => temp(12179 DOWNTO 12170) := ADC(11 DOWNTO 2);
			WHEN 1218 => temp(12189 DOWNTO 12180) := ADC(11 DOWNTO 2);
			WHEN 1219 => temp(12199 DOWNTO 12190) := ADC(11 DOWNTO 2);
			WHEN 1220 => temp(12209 DOWNTO 12200) := ADC(11 DOWNTO 2);
			WHEN 1221 => temp(12219 DOWNTO 12210) := ADC(11 DOWNTO 2);
			WHEN 1222 => temp(12229 DOWNTO 12220) := ADC(11 DOWNTO 2);
			WHEN 1223 => temp(12239 DOWNTO 12230) := ADC(11 DOWNTO 2);
			WHEN 1224 => temp(12249 DOWNTO 12240) := ADC(11 DOWNTO 2);
			WHEN 1225 => temp(12259 DOWNTO 12250) := ADC(11 DOWNTO 2);
			WHEN 1226 => temp(12269 DOWNTO 12260) := ADC(11 DOWNTO 2);
			WHEN 1227 => temp(12279 DOWNTO 12270) := ADC(11 DOWNTO 2);
			WHEN 1228 => temp(12289 DOWNTO 12280) := ADC(11 DOWNTO 2);
			WHEN 1229 => temp(12299 DOWNTO 12290) := ADC(11 DOWNTO 2);
			WHEN 1230 => temp(12309 DOWNTO 12300) := ADC(11 DOWNTO 2);
			WHEN 1231 => temp(12319 DOWNTO 12310) := ADC(11 DOWNTO 2);
			WHEN 1232 => temp(12329 DOWNTO 12320) := ADC(11 DOWNTO 2);
			WHEN 1233 => temp(12339 DOWNTO 12330) := ADC(11 DOWNTO 2);
			WHEN 1234 => temp(12349 DOWNTO 12340) := ADC(11 DOWNTO 2);
			WHEN 1235 => temp(12359 DOWNTO 12350) := ADC(11 DOWNTO 2);
			WHEN 1236 => temp(12369 DOWNTO 12360) := ADC(11 DOWNTO 2);
			WHEN 1237 => temp(12379 DOWNTO 12370) := ADC(11 DOWNTO 2);
			WHEN 1238 => temp(12389 DOWNTO 12380) := ADC(11 DOWNTO 2);
			WHEN 1239 => temp(12399 DOWNTO 12390) := ADC(11 DOWNTO 2);
			WHEN 1240 => temp(12409 DOWNTO 12400) := ADC(11 DOWNTO 2);
			WHEN 1241 => temp(12419 DOWNTO 12410) := ADC(11 DOWNTO 2);
			WHEN 1242 => temp(12429 DOWNTO 12420) := ADC(11 DOWNTO 2);
			WHEN 1243 => temp(12439 DOWNTO 12430) := ADC(11 DOWNTO 2);
			WHEN 1244 => temp(12449 DOWNTO 12440) := ADC(11 DOWNTO 2);
			WHEN 1245 => temp(12459 DOWNTO 12450) := ADC(11 DOWNTO 2);
			WHEN 1246 => temp(12469 DOWNTO 12460) := ADC(11 DOWNTO 2);
			WHEN 1247 => temp(12479 DOWNTO 12470) := ADC(11 DOWNTO 2);
			WHEN 1248 => temp(12489 DOWNTO 12480) := ADC(11 DOWNTO 2);
			WHEN 1249 => temp(12499 DOWNTO 12490) := ADC(11 DOWNTO 2);
			WHEN 1250 => temp(12509 DOWNTO 12500) := ADC(11 DOWNTO 2);
			WHEN 1251 => temp(12519 DOWNTO 12510) := ADC(11 DOWNTO 2);
			WHEN 1252 => temp(12529 DOWNTO 12520) := ADC(11 DOWNTO 2);
			WHEN 1253 => temp(12539 DOWNTO 12530) := ADC(11 DOWNTO 2);
			WHEN 1254 => temp(12549 DOWNTO 12540) := ADC(11 DOWNTO 2);
			WHEN 1255 => temp(12559 DOWNTO 12550) := ADC(11 DOWNTO 2);
			WHEN 1256 => temp(12569 DOWNTO 12560) := ADC(11 DOWNTO 2);
			WHEN 1257 => temp(12579 DOWNTO 12570) := ADC(11 DOWNTO 2);
			WHEN 1258 => temp(12589 DOWNTO 12580) := ADC(11 DOWNTO 2);
			WHEN 1259 => temp(12599 DOWNTO 12590) := ADC(11 DOWNTO 2);
			WHEN 1260 => temp(12609 DOWNTO 12600) := ADC(11 DOWNTO 2);
			WHEN 1261 => temp(12619 DOWNTO 12610) := ADC(11 DOWNTO 2);
			WHEN 1262 => temp(12629 DOWNTO 12620) := ADC(11 DOWNTO 2);
			WHEN 1263 => temp(12639 DOWNTO 12630) := ADC(11 DOWNTO 2);
			WHEN 1264 => temp(12649 DOWNTO 12640) := ADC(11 DOWNTO 2);
			WHEN 1265 => temp(12659 DOWNTO 12650) := ADC(11 DOWNTO 2);
			WHEN 1266 => temp(12669 DOWNTO 12660) := ADC(11 DOWNTO 2);
			WHEN 1267 => temp(12679 DOWNTO 12670) := ADC(11 DOWNTO 2);
			WHEN 1268 => temp(12689 DOWNTO 12680) := ADC(11 DOWNTO 2);
			WHEN 1269 => temp(12699 DOWNTO 12690) := ADC(11 DOWNTO 2);
			WHEN 1270 => temp(12709 DOWNTO 12700) := ADC(11 DOWNTO 2);
			WHEN 1271 => temp(12719 DOWNTO 12710) := ADC(11 DOWNTO 2);
			WHEN 1272 => temp(12729 DOWNTO 12720) := ADC(11 DOWNTO 2);
			WHEN 1273 => temp(12739 DOWNTO 12730) := ADC(11 DOWNTO 2);
			WHEN 1274 => temp(12749 DOWNTO 12740) := ADC(11 DOWNTO 2);
			WHEN 1275 => temp(12759 DOWNTO 12750) := ADC(11 DOWNTO 2);
			WHEN 1276 => temp(12769 DOWNTO 12760) := ADC(11 DOWNTO 2);
			WHEN 1277 => temp(12779 DOWNTO 12770) := ADC(11 DOWNTO 2);
			WHEN 1278 => temp(12789 DOWNTO 12780) := ADC(11 DOWNTO 2);
			WHEN 1279 => temp(12799 DOWNTO 12790) := ADC(11 DOWNTO 2);
			WHEN 1280 => temp(12809 DOWNTO 12800) := ADC(11 DOWNTO 2);
			WHEN 1281 => temp(12819 DOWNTO 12810) := ADC(11 DOWNTO 2);
			WHEN 1282 => temp(12829 DOWNTO 12820) := ADC(11 DOWNTO 2);
			WHEN 1283 => temp(12839 DOWNTO 12830) := ADC(11 DOWNTO 2);
			WHEN 1284 => temp(12849 DOWNTO 12840) := ADC(11 DOWNTO 2);
			WHEN 1285 => temp(12859 DOWNTO 12850) := ADC(11 DOWNTO 2);
			WHEN 1286 => temp(12869 DOWNTO 12860) := ADC(11 DOWNTO 2);
			WHEN 1287 => temp(12879 DOWNTO 12870) := ADC(11 DOWNTO 2);
			WHEN 1288 => temp(12889 DOWNTO 12880) := ADC(11 DOWNTO 2);
			WHEN 1289 => temp(12899 DOWNTO 12890) := ADC(11 DOWNTO 2);
			WHEN 1290 => temp(12909 DOWNTO 12900) := ADC(11 DOWNTO 2);
			WHEN 1291 => temp(12919 DOWNTO 12910) := ADC(11 DOWNTO 2);
			WHEN 1292 => temp(12929 DOWNTO 12920) := ADC(11 DOWNTO 2);
			WHEN 1293 => temp(12939 DOWNTO 12930) := ADC(11 DOWNTO 2);
			WHEN 1294 => temp(12949 DOWNTO 12940) := ADC(11 DOWNTO 2);
			WHEN 1295 => temp(12959 DOWNTO 12950) := ADC(11 DOWNTO 2);
			WHEN 1296 => temp(12969 DOWNTO 12960) := ADC(11 DOWNTO 2);
			WHEN 1297 => temp(12979 DOWNTO 12970) := ADC(11 DOWNTO 2);
			WHEN 1298 => temp(12989 DOWNTO 12980) := ADC(11 DOWNTO 2);
			WHEN 1299 => temp(12999 DOWNTO 12990) := ADC(11 DOWNTO 2);
			WHEN 1300 => temp(13009 DOWNTO 13000) := ADC(11 DOWNTO 2);
			WHEN 1301 => temp(13019 DOWNTO 13010) := ADC(11 DOWNTO 2);
			WHEN 1302 => temp(13029 DOWNTO 13020) := ADC(11 DOWNTO 2);
			WHEN 1303 => temp(13039 DOWNTO 13030) := ADC(11 DOWNTO 2);
			WHEN 1304 => temp(13049 DOWNTO 13040) := ADC(11 DOWNTO 2);
			WHEN 1305 => temp(13059 DOWNTO 13050) := ADC(11 DOWNTO 2);
			WHEN 1306 => temp(13069 DOWNTO 13060) := ADC(11 DOWNTO 2);
			WHEN 1307 => temp(13079 DOWNTO 13070) := ADC(11 DOWNTO 2);
			WHEN 1308 => temp(13089 DOWNTO 13080) := ADC(11 DOWNTO 2);
			WHEN 1309 => temp(13099 DOWNTO 13090) := ADC(11 DOWNTO 2);
			WHEN 1310 => temp(13109 DOWNTO 13100) := ADC(11 DOWNTO 2);
			WHEN 1311 => temp(13119 DOWNTO 13110) := ADC(11 DOWNTO 2);
			WHEN 1312 => temp(13129 DOWNTO 13120) := ADC(11 DOWNTO 2);
			WHEN 1313 => temp(13139 DOWNTO 13130) := ADC(11 DOWNTO 2);
			WHEN 1314 => temp(13149 DOWNTO 13140) := ADC(11 DOWNTO 2);
			WHEN 1315 => temp(13159 DOWNTO 13150) := ADC(11 DOWNTO 2);
			WHEN 1316 => temp(13169 DOWNTO 13160) := ADC(11 DOWNTO 2);
			WHEN 1317 => temp(13179 DOWNTO 13170) := ADC(11 DOWNTO 2);
			WHEN 1318 => temp(13189 DOWNTO 13180) := ADC(11 DOWNTO 2);
			WHEN 1319 => temp(13199 DOWNTO 13190) := ADC(11 DOWNTO 2);
			WHEN 1320 => temp(13209 DOWNTO 13200) := ADC(11 DOWNTO 2);
			WHEN 1321 => temp(13219 DOWNTO 13210) := ADC(11 DOWNTO 2);
			WHEN 1322 => temp(13229 DOWNTO 13220) := ADC(11 DOWNTO 2);
			WHEN 1323 => temp(13239 DOWNTO 13230) := ADC(11 DOWNTO 2);
			WHEN 1324 => temp(13249 DOWNTO 13240) := ADC(11 DOWNTO 2);
			WHEN 1325 => temp(13259 DOWNTO 13250) := ADC(11 DOWNTO 2);
			WHEN 1326 => temp(13269 DOWNTO 13260) := ADC(11 DOWNTO 2);
			WHEN 1327 => temp(13279 DOWNTO 13270) := ADC(11 DOWNTO 2);
			WHEN 1328 => temp(13289 DOWNTO 13280) := ADC(11 DOWNTO 2);
			WHEN 1329 => temp(13299 DOWNTO 13290) := ADC(11 DOWNTO 2);
			WHEN 1330 => temp(13309 DOWNTO 13300) := ADC(11 DOWNTO 2);
			WHEN 1331 => temp(13319 DOWNTO 13310) := ADC(11 DOWNTO 2);
			WHEN 1332 => temp(13329 DOWNTO 13320) := ADC(11 DOWNTO 2);
			WHEN 1333 => temp(13339 DOWNTO 13330) := ADC(11 DOWNTO 2);
			WHEN 1334 => temp(13349 DOWNTO 13340) := ADC(11 DOWNTO 2);
			WHEN 1335 => temp(13359 DOWNTO 13350) := ADC(11 DOWNTO 2);
			WHEN 1336 => temp(13369 DOWNTO 13360) := ADC(11 DOWNTO 2);
			WHEN 1337 => temp(13379 DOWNTO 13370) := ADC(11 DOWNTO 2);
			WHEN 1338 => temp(13389 DOWNTO 13380) := ADC(11 DOWNTO 2);
			WHEN 1339 => temp(13399 DOWNTO 13390) := ADC(11 DOWNTO 2);
			WHEN 1340 => temp(13409 DOWNTO 13400) := ADC(11 DOWNTO 2);
			WHEN 1341 => temp(13419 DOWNTO 13410) := ADC(11 DOWNTO 2);
			WHEN 1342 => temp(13429 DOWNTO 13420) := ADC(11 DOWNTO 2);
			WHEN 1343 => temp(13439 DOWNTO 13430) := ADC(11 DOWNTO 2);
			WHEN 1344 => temp(13449 DOWNTO 13440) := ADC(11 DOWNTO 2);
			WHEN 1345 => temp(13459 DOWNTO 13450) := ADC(11 DOWNTO 2);
			WHEN 1346 => temp(13469 DOWNTO 13460) := ADC(11 DOWNTO 2);
			WHEN 1347 => temp(13479 DOWNTO 13470) := ADC(11 DOWNTO 2);
			WHEN 1348 => temp(13489 DOWNTO 13480) := ADC(11 DOWNTO 2);
			WHEN 1349 => temp(13499 DOWNTO 13490) := ADC(11 DOWNTO 2);
			WHEN 1350 => temp(13509 DOWNTO 13500) := ADC(11 DOWNTO 2);
			WHEN 1351 => temp(13519 DOWNTO 13510) := ADC(11 DOWNTO 2);
			WHEN 1352 => temp(13529 DOWNTO 13520) := ADC(11 DOWNTO 2);
			WHEN 1353 => temp(13539 DOWNTO 13530) := ADC(11 DOWNTO 2);
			WHEN 1354 => temp(13549 DOWNTO 13540) := ADC(11 DOWNTO 2);
			WHEN 1355 => temp(13559 DOWNTO 13550) := ADC(11 DOWNTO 2);
			WHEN 1356 => temp(13569 DOWNTO 13560) := ADC(11 DOWNTO 2);
			WHEN 1357 => temp(13579 DOWNTO 13570) := ADC(11 DOWNTO 2);
			WHEN 1358 => temp(13589 DOWNTO 13580) := ADC(11 DOWNTO 2);
			WHEN 1359 => temp(13599 DOWNTO 13590) := ADC(11 DOWNTO 2);
			WHEN 1360 => temp(13609 DOWNTO 13600) := ADC(11 DOWNTO 2);
			WHEN 1361 => temp(13619 DOWNTO 13610) := ADC(11 DOWNTO 2);
			WHEN 1362 => temp(13629 DOWNTO 13620) := ADC(11 DOWNTO 2);
			WHEN 1363 => temp(13639 DOWNTO 13630) := ADC(11 DOWNTO 2);
			WHEN 1364 => temp(13649 DOWNTO 13640) := ADC(11 DOWNTO 2);
			WHEN 1365 => temp(13659 DOWNTO 13650) := ADC(11 DOWNTO 2);
			WHEN 1366 => temp(13669 DOWNTO 13660) := ADC(11 DOWNTO 2);
			WHEN 1367 => temp(13679 DOWNTO 13670) := ADC(11 DOWNTO 2);
			WHEN 1368 => temp(13689 DOWNTO 13680) := ADC(11 DOWNTO 2);
			WHEN 1369 => temp(13699 DOWNTO 13690) := ADC(11 DOWNTO 2);
			WHEN 1370 => temp(13709 DOWNTO 13700) := ADC(11 DOWNTO 2);
			WHEN 1371 => temp(13719 DOWNTO 13710) := ADC(11 DOWNTO 2);
			WHEN 1372 => temp(13729 DOWNTO 13720) := ADC(11 DOWNTO 2);
			WHEN 1373 => temp(13739 DOWNTO 13730) := ADC(11 DOWNTO 2);
			WHEN 1374 => temp(13749 DOWNTO 13740) := ADC(11 DOWNTO 2);
			WHEN 1375 => temp(13759 DOWNTO 13750) := ADC(11 DOWNTO 2);
			WHEN 1376 => temp(13769 DOWNTO 13760) := ADC(11 DOWNTO 2);
			WHEN 1377 => temp(13779 DOWNTO 13770) := ADC(11 DOWNTO 2);
			WHEN 1378 => temp(13789 DOWNTO 13780) := ADC(11 DOWNTO 2);
			WHEN 1379 => temp(13799 DOWNTO 13790) := ADC(11 DOWNTO 2);
			WHEN 1380 => temp(13809 DOWNTO 13800) := ADC(11 DOWNTO 2);
			WHEN 1381 => temp(13819 DOWNTO 13810) := ADC(11 DOWNTO 2);
			WHEN 1382 => temp(13829 DOWNTO 13820) := ADC(11 DOWNTO 2);
			WHEN 1383 => temp(13839 DOWNTO 13830) := ADC(11 DOWNTO 2);
			WHEN 1384 => temp(13849 DOWNTO 13840) := ADC(11 DOWNTO 2);
			WHEN 1385 => temp(13859 DOWNTO 13850) := ADC(11 DOWNTO 2);
			WHEN 1386 => temp(13869 DOWNTO 13860) := ADC(11 DOWNTO 2);
			WHEN 1387 => temp(13879 DOWNTO 13870) := ADC(11 DOWNTO 2);
			WHEN 1388 => temp(13889 DOWNTO 13880) := ADC(11 DOWNTO 2);
			WHEN 1389 => temp(13899 DOWNTO 13890) := ADC(11 DOWNTO 2);
			WHEN 1390 => temp(13909 DOWNTO 13900) := ADC(11 DOWNTO 2);
			WHEN 1391 => temp(13919 DOWNTO 13910) := ADC(11 DOWNTO 2);
			WHEN 1392 => temp(13929 DOWNTO 13920) := ADC(11 DOWNTO 2);
			WHEN 1393 => temp(13939 DOWNTO 13930) := ADC(11 DOWNTO 2);
			WHEN 1394 => temp(13949 DOWNTO 13940) := ADC(11 DOWNTO 2);
			WHEN 1395 => temp(13959 DOWNTO 13950) := ADC(11 DOWNTO 2);
			WHEN 1396 => temp(13969 DOWNTO 13960) := ADC(11 DOWNTO 2);
			WHEN 1397 => temp(13979 DOWNTO 13970) := ADC(11 DOWNTO 2);
			WHEN 1398 => temp(13989 DOWNTO 13980) := ADC(11 DOWNTO 2);
			WHEN 1399 => temp(13999 DOWNTO 13990) := ADC(11 DOWNTO 2);
			WHEN 1400 => temp(14009 DOWNTO 14000) := ADC(11 DOWNTO 2);
			WHEN 1401 => temp(14019 DOWNTO 14010) := ADC(11 DOWNTO 2);
			WHEN 1402 => temp(14029 DOWNTO 14020) := ADC(11 DOWNTO 2);
			WHEN 1403 => temp(14039 DOWNTO 14030) := ADC(11 DOWNTO 2);
			WHEN 1404 => temp(14049 DOWNTO 14040) := ADC(11 DOWNTO 2);
			WHEN 1405 => temp(14059 DOWNTO 14050) := ADC(11 DOWNTO 2);
			WHEN 1406 => temp(14069 DOWNTO 14060) := ADC(11 DOWNTO 2);
			WHEN 1407 => temp(14079 DOWNTO 14070) := ADC(11 DOWNTO 2);
			WHEN 1408 => temp(14089 DOWNTO 14080) := ADC(11 DOWNTO 2);
			WHEN 1409 => temp(14099 DOWNTO 14090) := ADC(11 DOWNTO 2);
			WHEN 1410 => temp(14109 DOWNTO 14100) := ADC(11 DOWNTO 2);
			WHEN 1411 => temp(14119 DOWNTO 14110) := ADC(11 DOWNTO 2);
			WHEN 1412 => temp(14129 DOWNTO 14120) := ADC(11 DOWNTO 2);
			WHEN 1413 => temp(14139 DOWNTO 14130) := ADC(11 DOWNTO 2);
			WHEN 1414 => temp(14149 DOWNTO 14140) := ADC(11 DOWNTO 2);
			WHEN 1415 => temp(14159 DOWNTO 14150) := ADC(11 DOWNTO 2);
			WHEN 1416 => temp(14169 DOWNTO 14160) := ADC(11 DOWNTO 2);
			WHEN 1417 => temp(14179 DOWNTO 14170) := ADC(11 DOWNTO 2);
			WHEN 1418 => temp(14189 DOWNTO 14180) := ADC(11 DOWNTO 2);
			WHEN 1419 => temp(14199 DOWNTO 14190) := ADC(11 DOWNTO 2);
			WHEN 1420 => temp(14209 DOWNTO 14200) := ADC(11 DOWNTO 2);
			WHEN 1421 => temp(14219 DOWNTO 14210) := ADC(11 DOWNTO 2);
			WHEN 1422 => temp(14229 DOWNTO 14220) := ADC(11 DOWNTO 2);
			WHEN 1423 => temp(14239 DOWNTO 14230) := ADC(11 DOWNTO 2);
			WHEN 1424 => temp(14249 DOWNTO 14240) := ADC(11 DOWNTO 2);
			WHEN 1425 => temp(14259 DOWNTO 14250) := ADC(11 DOWNTO 2);
			WHEN 1426 => temp(14269 DOWNTO 14260) := ADC(11 DOWNTO 2);
			WHEN 1427 => temp(14279 DOWNTO 14270) := ADC(11 DOWNTO 2);
			WHEN 1428 => temp(14289 DOWNTO 14280) := ADC(11 DOWNTO 2);
			WHEN 1429 => temp(14299 DOWNTO 14290) := ADC(11 DOWNTO 2);
			WHEN 1430 => temp(14309 DOWNTO 14300) := ADC(11 DOWNTO 2);
			WHEN 1431 => temp(14319 DOWNTO 14310) := ADC(11 DOWNTO 2);
			WHEN 1432 => temp(14329 DOWNTO 14320) := ADC(11 DOWNTO 2);
			WHEN 1433 => temp(14339 DOWNTO 14330) := ADC(11 DOWNTO 2);
			WHEN 1434 => temp(14349 DOWNTO 14340) := ADC(11 DOWNTO 2);
			WHEN 1435 => temp(14359 DOWNTO 14350) := ADC(11 DOWNTO 2);
			WHEN 1436 => temp(14369 DOWNTO 14360) := ADC(11 DOWNTO 2);
			WHEN 1437 => temp(14379 DOWNTO 14370) := ADC(11 DOWNTO 2);
			WHEN 1438 => temp(14389 DOWNTO 14380) := ADC(11 DOWNTO 2);
			WHEN 1439 => temp(14399 DOWNTO 14390) := ADC(11 DOWNTO 2);
			WHEN 1440 => temp(14409 DOWNTO 14400) := ADC(11 DOWNTO 2);
			WHEN 1441 => temp(14419 DOWNTO 14410) := ADC(11 DOWNTO 2);
			WHEN 1442 => temp(14429 DOWNTO 14420) := ADC(11 DOWNTO 2);
			WHEN 1443 => temp(14439 DOWNTO 14430) := ADC(11 DOWNTO 2);
			WHEN 1444 => temp(14449 DOWNTO 14440) := ADC(11 DOWNTO 2);
			WHEN 1445 => temp(14459 DOWNTO 14450) := ADC(11 DOWNTO 2);
			WHEN 1446 => temp(14469 DOWNTO 14460) := ADC(11 DOWNTO 2);
			WHEN 1447 => temp(14479 DOWNTO 14470) := ADC(11 DOWNTO 2);
			WHEN 1448 => temp(14489 DOWNTO 14480) := ADC(11 DOWNTO 2);
			WHEN 1449 => temp(14499 DOWNTO 14490) := ADC(11 DOWNTO 2);
			WHEN 1450 => temp(14509 DOWNTO 14500) := ADC(11 DOWNTO 2);
			WHEN 1451 => temp(14519 DOWNTO 14510) := ADC(11 DOWNTO 2);
			WHEN 1452 => temp(14529 DOWNTO 14520) := ADC(11 DOWNTO 2);
			WHEN 1453 => temp(14539 DOWNTO 14530) := ADC(11 DOWNTO 2);
			WHEN 1454 => temp(14549 DOWNTO 14540) := ADC(11 DOWNTO 2);
			WHEN 1455 => temp(14559 DOWNTO 14550) := ADC(11 DOWNTO 2);
			WHEN 1456 => temp(14569 DOWNTO 14560) := ADC(11 DOWNTO 2);
			WHEN 1457 => temp(14579 DOWNTO 14570) := ADC(11 DOWNTO 2);
			WHEN 1458 => temp(14589 DOWNTO 14580) := ADC(11 DOWNTO 2);
			WHEN 1459 => temp(14599 DOWNTO 14590) := ADC(11 DOWNTO 2);
			WHEN 1460 => temp(14609 DOWNTO 14600) := ADC(11 DOWNTO 2);
			WHEN 1461 => temp(14619 DOWNTO 14610) := ADC(11 DOWNTO 2);
			WHEN 1462 => temp(14629 DOWNTO 14620) := ADC(11 DOWNTO 2);
			WHEN 1463 => temp(14639 DOWNTO 14630) := ADC(11 DOWNTO 2);
			WHEN 1464 => temp(14649 DOWNTO 14640) := ADC(11 DOWNTO 2);
			WHEN 1465 => temp(14659 DOWNTO 14650) := ADC(11 DOWNTO 2);
			WHEN 1466 => temp(14669 DOWNTO 14660) := ADC(11 DOWNTO 2);
			WHEN 1467 => temp(14679 DOWNTO 14670) := ADC(11 DOWNTO 2);
			WHEN 1468 => temp(14689 DOWNTO 14680) := ADC(11 DOWNTO 2);
			WHEN 1469 => temp(14699 DOWNTO 14690) := ADC(11 DOWNTO 2);
			WHEN 1470 => temp(14709 DOWNTO 14700) := ADC(11 DOWNTO 2);
			WHEN 1471 => temp(14719 DOWNTO 14710) := ADC(11 DOWNTO 2);
			WHEN 1472 => temp(14729 DOWNTO 14720) := ADC(11 DOWNTO 2);
			WHEN 1473 => temp(14739 DOWNTO 14730) := ADC(11 DOWNTO 2);
			WHEN 1474 => temp(14749 DOWNTO 14740) := ADC(11 DOWNTO 2);
			WHEN 1475 => temp(14759 DOWNTO 14750) := ADC(11 DOWNTO 2);
			WHEN 1476 => temp(14769 DOWNTO 14760) := ADC(11 DOWNTO 2);
			WHEN 1477 => temp(14779 DOWNTO 14770) := ADC(11 DOWNTO 2);
			WHEN 1478 => temp(14789 DOWNTO 14780) := ADC(11 DOWNTO 2);
			WHEN 1479 => temp(14799 DOWNTO 14790) := ADC(11 DOWNTO 2);
			WHEN 1480 => temp(14809 DOWNTO 14800) := ADC(11 DOWNTO 2);
			WHEN 1481 => temp(14819 DOWNTO 14810) := ADC(11 DOWNTO 2);
			WHEN 1482 => temp(14829 DOWNTO 14820) := ADC(11 DOWNTO 2);
			WHEN 1483 => temp(14839 DOWNTO 14830) := ADC(11 DOWNTO 2);
			WHEN 1484 => temp(14849 DOWNTO 14840) := ADC(11 DOWNTO 2);
			WHEN 1485 => temp(14859 DOWNTO 14850) := ADC(11 DOWNTO 2);
			WHEN 1486 => temp(14869 DOWNTO 14860) := ADC(11 DOWNTO 2);
			WHEN 1487 => temp(14879 DOWNTO 14870) := ADC(11 DOWNTO 2);
			WHEN 1488 => temp(14889 DOWNTO 14880) := ADC(11 DOWNTO 2);
			WHEN 1489 => temp(14899 DOWNTO 14890) := ADC(11 DOWNTO 2);
			WHEN 1490 => temp(14909 DOWNTO 14900) := ADC(11 DOWNTO 2);
			WHEN 1491 => temp(14919 DOWNTO 14910) := ADC(11 DOWNTO 2);
			WHEN 1492 => temp(14929 DOWNTO 14920) := ADC(11 DOWNTO 2);
			WHEN 1493 => temp(14939 DOWNTO 14930) := ADC(11 DOWNTO 2);
			WHEN 1494 => temp(14949 DOWNTO 14940) := ADC(11 DOWNTO 2);
			WHEN 1495 => temp(14959 DOWNTO 14950) := ADC(11 DOWNTO 2);
			WHEN 1496 => temp(14969 DOWNTO 14960) := ADC(11 DOWNTO 2);
			WHEN 1497 => temp(14979 DOWNTO 14970) := ADC(11 DOWNTO 2);
			WHEN 1498 => temp(14989 DOWNTO 14980) := ADC(11 DOWNTO 2);
			WHEN 1499 => temp(14999 DOWNTO 14990) := ADC(11 DOWNTO 2);
			WHEN 1500 => temp(15009 DOWNTO 15000) := ADC(11 DOWNTO 2);
			WHEN 1501 => temp(15019 DOWNTO 15010) := ADC(11 DOWNTO 2);
			WHEN 1502 => temp(15029 DOWNTO 15020) := ADC(11 DOWNTO 2);
			WHEN 1503 => temp(15039 DOWNTO 15030) := ADC(11 DOWNTO 2);
			WHEN 1504 => temp(15049 DOWNTO 15040) := ADC(11 DOWNTO 2);
			WHEN 1505 => temp(15059 DOWNTO 15050) := ADC(11 DOWNTO 2);
			WHEN 1506 => temp(15069 DOWNTO 15060) := ADC(11 DOWNTO 2);
			WHEN 1507 => temp(15079 DOWNTO 15070) := ADC(11 DOWNTO 2);
			WHEN 1508 => temp(15089 DOWNTO 15080) := ADC(11 DOWNTO 2);
			WHEN 1509 => temp(15099 DOWNTO 15090) := ADC(11 DOWNTO 2);
			WHEN 1510 => temp(15109 DOWNTO 15100) := ADC(11 DOWNTO 2);
			WHEN 1511 => temp(15119 DOWNTO 15110) := ADC(11 DOWNTO 2);
			WHEN 1512 => temp(15129 DOWNTO 15120) := ADC(11 DOWNTO 2);
			WHEN 1513 => temp(15139 DOWNTO 15130) := ADC(11 DOWNTO 2);
			WHEN 1514 => temp(15149 DOWNTO 15140) := ADC(11 DOWNTO 2);
			WHEN 1515 => temp(15159 DOWNTO 15150) := ADC(11 DOWNTO 2);
			WHEN 1516 => temp(15169 DOWNTO 15160) := ADC(11 DOWNTO 2);
			WHEN 1517 => temp(15179 DOWNTO 15170) := ADC(11 DOWNTO 2);
			WHEN 1518 => temp(15189 DOWNTO 15180) := ADC(11 DOWNTO 2);
			WHEN 1519 => temp(15199 DOWNTO 15190) := ADC(11 DOWNTO 2);
			WHEN 1520 => temp(15209 DOWNTO 15200) := ADC(11 DOWNTO 2);
			WHEN 1521 => temp(15219 DOWNTO 15210) := ADC(11 DOWNTO 2);
			WHEN 1522 => temp(15229 DOWNTO 15220) := ADC(11 DOWNTO 2);
			WHEN 1523 => temp(15239 DOWNTO 15230) := ADC(11 DOWNTO 2);
			WHEN 1524 => temp(15249 DOWNTO 15240) := ADC(11 DOWNTO 2);
			WHEN 1525 => temp(15259 DOWNTO 15250) := ADC(11 DOWNTO 2);
			WHEN 1526 => temp(15269 DOWNTO 15260) := ADC(11 DOWNTO 2);
			WHEN 1527 => temp(15279 DOWNTO 15270) := ADC(11 DOWNTO 2);
			WHEN 1528 => temp(15289 DOWNTO 15280) := ADC(11 DOWNTO 2);
			WHEN 1529 => temp(15299 DOWNTO 15290) := ADC(11 DOWNTO 2);
			WHEN 1530 => temp(15309 DOWNTO 15300) := ADC(11 DOWNTO 2);
			WHEN 1531 => temp(15319 DOWNTO 15310) := ADC(11 DOWNTO 2);
			WHEN 1532 => temp(15329 DOWNTO 15320) := ADC(11 DOWNTO 2);
			WHEN 1533 => temp(15339 DOWNTO 15330) := ADC(11 DOWNTO 2);
			WHEN 1534 => temp(15349 DOWNTO 15340) := ADC(11 DOWNTO 2);
			WHEN 1535 => temp(15359 DOWNTO 15350) := ADC(11 DOWNTO 2);
			WHEN 1536 => temp(15369 DOWNTO 15360) := ADC(11 DOWNTO 2);
			WHEN 1537 => temp(15379 DOWNTO 15370) := ADC(11 DOWNTO 2);
			WHEN 1538 => temp(15389 DOWNTO 15380) := ADC(11 DOWNTO 2);
			WHEN 1539 => temp(15399 DOWNTO 15390) := ADC(11 DOWNTO 2);
			WHEN 1540 => temp(15409 DOWNTO 15400) := ADC(11 DOWNTO 2);
			WHEN 1541 => temp(15419 DOWNTO 15410) := ADC(11 DOWNTO 2);
			WHEN 1542 => temp(15429 DOWNTO 15420) := ADC(11 DOWNTO 2);
			WHEN 1543 => temp(15439 DOWNTO 15430) := ADC(11 DOWNTO 2);
			WHEN 1544 => temp(15449 DOWNTO 15440) := ADC(11 DOWNTO 2);
			WHEN 1545 => temp(15459 DOWNTO 15450) := ADC(11 DOWNTO 2);
			WHEN 1546 => temp(15469 DOWNTO 15460) := ADC(11 DOWNTO 2);
			WHEN 1547 => temp(15479 DOWNTO 15470) := ADC(11 DOWNTO 2);
			WHEN 1548 => temp(15489 DOWNTO 15480) := ADC(11 DOWNTO 2);
			WHEN 1549 => temp(15499 DOWNTO 15490) := ADC(11 DOWNTO 2);
			WHEN 1550 => temp(15509 DOWNTO 15500) := ADC(11 DOWNTO 2);
			WHEN 1551 => temp(15519 DOWNTO 15510) := ADC(11 DOWNTO 2);
			WHEN 1552 => temp(15529 DOWNTO 15520) := ADC(11 DOWNTO 2);
			WHEN 1553 => temp(15539 DOWNTO 15530) := ADC(11 DOWNTO 2);
			WHEN 1554 => temp(15549 DOWNTO 15540) := ADC(11 DOWNTO 2);
			WHEN 1555 => temp(15559 DOWNTO 15550) := ADC(11 DOWNTO 2);
			WHEN 1556 => temp(15569 DOWNTO 15560) := ADC(11 DOWNTO 2);
			WHEN 1557 => temp(15579 DOWNTO 15570) := ADC(11 DOWNTO 2);
			WHEN 1558 => temp(15589 DOWNTO 15580) := ADC(11 DOWNTO 2);
			WHEN 1559 => temp(15599 DOWNTO 15590) := ADC(11 DOWNTO 2);
			WHEN 1560 => temp(15609 DOWNTO 15600) := ADC(11 DOWNTO 2);
			WHEN 1561 => temp(15619 DOWNTO 15610) := ADC(11 DOWNTO 2);
			WHEN 1562 => temp(15629 DOWNTO 15620) := ADC(11 DOWNTO 2);
			WHEN 1563 => temp(15639 DOWNTO 15630) := ADC(11 DOWNTO 2);
			WHEN 1564 => temp(15649 DOWNTO 15640) := ADC(11 DOWNTO 2);
			WHEN 1565 => temp(15659 DOWNTO 15650) := ADC(11 DOWNTO 2);
			WHEN 1566 => temp(15669 DOWNTO 15660) := ADC(11 DOWNTO 2);
			WHEN 1567 => temp(15679 DOWNTO 15670) := ADC(11 DOWNTO 2);
			WHEN 1568 => temp(15689 DOWNTO 15680) := ADC(11 DOWNTO 2);
			WHEN 1569 => temp(15699 DOWNTO 15690) := ADC(11 DOWNTO 2);
			WHEN 1570 => temp(15709 DOWNTO 15700) := ADC(11 DOWNTO 2);
			WHEN 1571 => temp(15719 DOWNTO 15710) := ADC(11 DOWNTO 2);
			WHEN 1572 => temp(15729 DOWNTO 15720) := ADC(11 DOWNTO 2);
			WHEN 1573 => temp(15739 DOWNTO 15730) := ADC(11 DOWNTO 2);
			WHEN 1574 => temp(15749 DOWNTO 15740) := ADC(11 DOWNTO 2);
			WHEN 1575 => temp(15759 DOWNTO 15750) := ADC(11 DOWNTO 2);
			WHEN 1576 => temp(15769 DOWNTO 15760) := ADC(11 DOWNTO 2);
			WHEN 1577 => temp(15779 DOWNTO 15770) := ADC(11 DOWNTO 2);
			WHEN 1578 => temp(15789 DOWNTO 15780) := ADC(11 DOWNTO 2);
			WHEN 1579 => temp(15799 DOWNTO 15790) := ADC(11 DOWNTO 2);
			WHEN 1580 => temp(15809 DOWNTO 15800) := ADC(11 DOWNTO 2);
			WHEN 1581 => temp(15819 DOWNTO 15810) := ADC(11 DOWNTO 2);
			WHEN 1582 => temp(15829 DOWNTO 15820) := ADC(11 DOWNTO 2);
			WHEN 1583 => temp(15839 DOWNTO 15830) := ADC(11 DOWNTO 2);
			WHEN 1584 => temp(15849 DOWNTO 15840) := ADC(11 DOWNTO 2);
			WHEN 1585 => temp(15859 DOWNTO 15850) := ADC(11 DOWNTO 2);
			WHEN 1586 => temp(15869 DOWNTO 15860) := ADC(11 DOWNTO 2);
			WHEN 1587 => temp(15879 DOWNTO 15870) := ADC(11 DOWNTO 2);
			WHEN 1588 => temp(15889 DOWNTO 15880) := ADC(11 DOWNTO 2);
			WHEN 1589 => temp(15899 DOWNTO 15890) := ADC(11 DOWNTO 2);
			WHEN 1590 => temp(15909 DOWNTO 15900) := ADC(11 DOWNTO 2);
			WHEN 1591 => temp(15919 DOWNTO 15910) := ADC(11 DOWNTO 2);
			WHEN 1592 => temp(15929 DOWNTO 15920) := ADC(11 DOWNTO 2);
			WHEN 1593 => temp(15939 DOWNTO 15930) := ADC(11 DOWNTO 2);
			WHEN 1594 => temp(15949 DOWNTO 15940) := ADC(11 DOWNTO 2);
			WHEN 1595 => temp(15959 DOWNTO 15950) := ADC(11 DOWNTO 2);
			WHEN 1596 => temp(15969 DOWNTO 15960) := ADC(11 DOWNTO 2);
			WHEN 1597 => temp(15979 DOWNTO 15970) := ADC(11 DOWNTO 2);
			WHEN 1598 => temp(15989 DOWNTO 15980) := ADC(11 DOWNTO 2);
			WHEN 1599 => temp(15999 DOWNTO 15990) := ADC(11 DOWNTO 2);
			WHEN 1600 => temp(16009 DOWNTO 16000) := ADC(11 DOWNTO 2);
			WHEN 1601 => temp(16019 DOWNTO 16010) := ADC(11 DOWNTO 2);
			WHEN 1602 => temp(16029 DOWNTO 16020) := ADC(11 DOWNTO 2);
			WHEN 1603 => temp(16039 DOWNTO 16030) := ADC(11 DOWNTO 2);
			WHEN 1604 => temp(16049 DOWNTO 16040) := ADC(11 DOWNTO 2);
			WHEN 1605 => temp(16059 DOWNTO 16050) := ADC(11 DOWNTO 2);
			WHEN 1606 => temp(16069 DOWNTO 16060) := ADC(11 DOWNTO 2);
			WHEN 1607 => temp(16079 DOWNTO 16070) := ADC(11 DOWNTO 2);
			WHEN 1608 => temp(16089 DOWNTO 16080) := ADC(11 DOWNTO 2);
			WHEN 1609 => temp(16099 DOWNTO 16090) := ADC(11 DOWNTO 2);
			WHEN 1610 => temp(16109 DOWNTO 16100) := ADC(11 DOWNTO 2);
			WHEN 1611 => temp(16119 DOWNTO 16110) := ADC(11 DOWNTO 2);
			WHEN 1612 => temp(16129 DOWNTO 16120) := ADC(11 DOWNTO 2);
			WHEN 1613 => temp(16139 DOWNTO 16130) := ADC(11 DOWNTO 2);
			WHEN 1614 => temp(16149 DOWNTO 16140) := ADC(11 DOWNTO 2);
			WHEN 1615 => temp(16159 DOWNTO 16150) := ADC(11 DOWNTO 2);
			WHEN 1616 => temp(16169 DOWNTO 16160) := ADC(11 DOWNTO 2);
			WHEN 1617 => temp(16179 DOWNTO 16170) := ADC(11 DOWNTO 2);
			WHEN 1618 => temp(16189 DOWNTO 16180) := ADC(11 DOWNTO 2);
			WHEN 1619 => temp(16199 DOWNTO 16190) := ADC(11 DOWNTO 2);
			WHEN 1620 => temp(16209 DOWNTO 16200) := ADC(11 DOWNTO 2);
			WHEN 1621 => temp(16219 DOWNTO 16210) := ADC(11 DOWNTO 2);
			WHEN 1622 => temp(16229 DOWNTO 16220) := ADC(11 DOWNTO 2);
			WHEN 1623 => temp(16239 DOWNTO 16230) := ADC(11 DOWNTO 2);
			WHEN 1624 => temp(16249 DOWNTO 16240) := ADC(11 DOWNTO 2);
			WHEN 1625 => temp(16259 DOWNTO 16250) := ADC(11 DOWNTO 2);
			WHEN 1626 => temp(16269 DOWNTO 16260) := ADC(11 DOWNTO 2);
			WHEN 1627 => temp(16279 DOWNTO 16270) := ADC(11 DOWNTO 2);
			WHEN 1628 => temp(16289 DOWNTO 16280) := ADC(11 DOWNTO 2);
			WHEN 1629 => temp(16299 DOWNTO 16290) := ADC(11 DOWNTO 2);
			WHEN 1630 => temp(16309 DOWNTO 16300) := ADC(11 DOWNTO 2);
			WHEN 1631 => temp(16319 DOWNTO 16310) := ADC(11 DOWNTO 2);
			WHEN 1632 => temp(16329 DOWNTO 16320) := ADC(11 DOWNTO 2);
			WHEN 1633 => temp(16339 DOWNTO 16330) := ADC(11 DOWNTO 2);
			WHEN 1634 => temp(16349 DOWNTO 16340) := ADC(11 DOWNTO 2);
			WHEN 1635 => temp(16359 DOWNTO 16350) := ADC(11 DOWNTO 2);
			WHEN 1636 => temp(16369 DOWNTO 16360) := ADC(11 DOWNTO 2);
			WHEN 1637 => temp(16379 DOWNTO 16370) := ADC(11 DOWNTO 2);
			WHEN 1638 => temp(16389 DOWNTO 16380) := ADC(11 DOWNTO 2);
			WHEN 1639 => temp(16399 DOWNTO 16390) := ADC(11 DOWNTO 2);
			WHEN 1640 => temp(16409 DOWNTO 16400) := ADC(11 DOWNTO 2);
			WHEN 1641 => temp(16419 DOWNTO 16410) := ADC(11 DOWNTO 2);
			WHEN 1642 => temp(16429 DOWNTO 16420) := ADC(11 DOWNTO 2);
			WHEN 1643 => temp(16439 DOWNTO 16430) := ADC(11 DOWNTO 2);
			WHEN 1644 => temp(16449 DOWNTO 16440) := ADC(11 DOWNTO 2);
			WHEN 1645 => temp(16459 DOWNTO 16450) := ADC(11 DOWNTO 2);
			WHEN 1646 => temp(16469 DOWNTO 16460) := ADC(11 DOWNTO 2);
			WHEN 1647 => temp(16479 DOWNTO 16470) := ADC(11 DOWNTO 2);
			WHEN 1648 => temp(16489 DOWNTO 16480) := ADC(11 DOWNTO 2);
			WHEN 1649 => temp(16499 DOWNTO 16490) := ADC(11 DOWNTO 2);
			WHEN 1650 => temp(16509 DOWNTO 16500) := ADC(11 DOWNTO 2);
			WHEN 1651 => temp(16519 DOWNTO 16510) := ADC(11 DOWNTO 2);
			WHEN 1652 => temp(16529 DOWNTO 16520) := ADC(11 DOWNTO 2);
			WHEN 1653 => temp(16539 DOWNTO 16530) := ADC(11 DOWNTO 2);
			WHEN 1654 => temp(16549 DOWNTO 16540) := ADC(11 DOWNTO 2);
			WHEN 1655 => temp(16559 DOWNTO 16550) := ADC(11 DOWNTO 2);
			WHEN 1656 => temp(16569 DOWNTO 16560) := ADC(11 DOWNTO 2);
			WHEN 1657 => temp(16579 DOWNTO 16570) := ADC(11 DOWNTO 2);
			WHEN 1658 => temp(16589 DOWNTO 16580) := ADC(11 DOWNTO 2);
			WHEN 1659 => temp(16599 DOWNTO 16590) := ADC(11 DOWNTO 2);
			WHEN 1660 => temp(16609 DOWNTO 16600) := ADC(11 DOWNTO 2);
			WHEN 1661 => temp(16619 DOWNTO 16610) := ADC(11 DOWNTO 2);
			WHEN 1662 => temp(16629 DOWNTO 16620) := ADC(11 DOWNTO 2);
			WHEN 1663 => temp(16639 DOWNTO 16630) := ADC(11 DOWNTO 2);
			WHEN 1664 => temp(16649 DOWNTO 16640) := ADC(11 DOWNTO 2);
			WHEN 1665 => temp(16659 DOWNTO 16650) := ADC(11 DOWNTO 2);
			WHEN 1666 => temp(16669 DOWNTO 16660) := ADC(11 DOWNTO 2);
			WHEN 1667 => temp(16679 DOWNTO 16670) := ADC(11 DOWNTO 2);
			WHEN 1668 => temp(16689 DOWNTO 16680) := ADC(11 DOWNTO 2);
			WHEN 1669 => temp(16699 DOWNTO 16690) := ADC(11 DOWNTO 2);
			WHEN 1670 => temp(16709 DOWNTO 16700) := ADC(11 DOWNTO 2);
			WHEN 1671 => temp(16719 DOWNTO 16710) := ADC(11 DOWNTO 2);
			WHEN 1672 => temp(16729 DOWNTO 16720) := ADC(11 DOWNTO 2);
			WHEN 1673 => temp(16739 DOWNTO 16730) := ADC(11 DOWNTO 2);
			WHEN 1674 => temp(16749 DOWNTO 16740) := ADC(11 DOWNTO 2);
			WHEN 1675 => temp(16759 DOWNTO 16750) := ADC(11 DOWNTO 2);
			WHEN 1676 => temp(16769 DOWNTO 16760) := ADC(11 DOWNTO 2);
			WHEN 1677 => temp(16779 DOWNTO 16770) := ADC(11 DOWNTO 2);
			WHEN 1678 => temp(16789 DOWNTO 16780) := ADC(11 DOWNTO 2);
			WHEN 1679 => temp(16799 DOWNTO 16790) := ADC(11 DOWNTO 2);
			WHEN 1680 => temp(16809 DOWNTO 16800) := ADC(11 DOWNTO 2);
			WHEN 1681 => temp(16819 DOWNTO 16810) := ADC(11 DOWNTO 2);
			WHEN 1682 => temp(16829 DOWNTO 16820) := ADC(11 DOWNTO 2);
			WHEN 1683 => temp(16839 DOWNTO 16830) := ADC(11 DOWNTO 2);
			WHEN 1684 => temp(16849 DOWNTO 16840) := ADC(11 DOWNTO 2);
			WHEN 1685 => temp(16859 DOWNTO 16850) := ADC(11 DOWNTO 2);
			WHEN 1686 => temp(16869 DOWNTO 16860) := ADC(11 DOWNTO 2);
			WHEN 1687 => temp(16879 DOWNTO 16870) := ADC(11 DOWNTO 2);
			WHEN 1688 => temp(16889 DOWNTO 16880) := ADC(11 DOWNTO 2);
			WHEN 1689 => temp(16899 DOWNTO 16890) := ADC(11 DOWNTO 2);
			WHEN 1690 => temp(16909 DOWNTO 16900) := ADC(11 DOWNTO 2);
			WHEN 1691 => temp(16919 DOWNTO 16910) := ADC(11 DOWNTO 2);
			WHEN 1692 => temp(16929 DOWNTO 16920) := ADC(11 DOWNTO 2);
			WHEN 1693 => temp(16939 DOWNTO 16930) := ADC(11 DOWNTO 2);
			WHEN 1694 => temp(16949 DOWNTO 16940) := ADC(11 DOWNTO 2);
			WHEN 1695 => temp(16959 DOWNTO 16950) := ADC(11 DOWNTO 2);
			WHEN 1696 => temp(16969 DOWNTO 16960) := ADC(11 DOWNTO 2);
			WHEN 1697 => temp(16979 DOWNTO 16970) := ADC(11 DOWNTO 2);
			WHEN 1698 => temp(16989 DOWNTO 16980) := ADC(11 DOWNTO 2);
			WHEN 1699 => temp(16999 DOWNTO 16990) := ADC(11 DOWNTO 2);
			WHEN 1700 => temp(17009 DOWNTO 17000) := ADC(11 DOWNTO 2);
			WHEN 1701 => temp(17019 DOWNTO 17010) := ADC(11 DOWNTO 2);
			WHEN 1702 => temp(17029 DOWNTO 17020) := ADC(11 DOWNTO 2);
			WHEN 1703 => temp(17039 DOWNTO 17030) := ADC(11 DOWNTO 2);
			WHEN 1704 => temp(17049 DOWNTO 17040) := ADC(11 DOWNTO 2);
			WHEN 1705 => temp(17059 DOWNTO 17050) := ADC(11 DOWNTO 2);
			WHEN 1706 => temp(17069 DOWNTO 17060) := ADC(11 DOWNTO 2);
			WHEN 1707 => temp(17079 DOWNTO 17070) := ADC(11 DOWNTO 2);
			WHEN 1708 => temp(17089 DOWNTO 17080) := ADC(11 DOWNTO 2);
			WHEN 1709 => temp(17099 DOWNTO 17090) := ADC(11 DOWNTO 2);
			WHEN 1710 => temp(17109 DOWNTO 17100) := ADC(11 DOWNTO 2);
			WHEN 1711 => temp(17119 DOWNTO 17110) := ADC(11 DOWNTO 2);
			WHEN 1712 => temp(17129 DOWNTO 17120) := ADC(11 DOWNTO 2);
			WHEN 1713 => temp(17139 DOWNTO 17130) := ADC(11 DOWNTO 2);
			WHEN 1714 => temp(17149 DOWNTO 17140) := ADC(11 DOWNTO 2);
			WHEN 1715 => temp(17159 DOWNTO 17150) := ADC(11 DOWNTO 2);
			WHEN 1716 => temp(17169 DOWNTO 17160) := ADC(11 DOWNTO 2);
			WHEN 1717 => temp(17179 DOWNTO 17170) := ADC(11 DOWNTO 2);
			WHEN 1718 => temp(17189 DOWNTO 17180) := ADC(11 DOWNTO 2);
			WHEN 1719 => temp(17199 DOWNTO 17190) := ADC(11 DOWNTO 2);
			WHEN 1720 => temp(17209 DOWNTO 17200) := ADC(11 DOWNTO 2);
			WHEN 1721 => temp(17219 DOWNTO 17210) := ADC(11 DOWNTO 2);
			WHEN 1722 => temp(17229 DOWNTO 17220) := ADC(11 DOWNTO 2);
			WHEN 1723 => temp(17239 DOWNTO 17230) := ADC(11 DOWNTO 2);
			WHEN 1724 => temp(17249 DOWNTO 17240) := ADC(11 DOWNTO 2);
			WHEN 1725 => temp(17259 DOWNTO 17250) := ADC(11 DOWNTO 2);
			WHEN 1726 => temp(17269 DOWNTO 17260) := ADC(11 DOWNTO 2);
			WHEN 1727 => temp(17279 DOWNTO 17270) := ADC(11 DOWNTO 2);
			WHEN 1728 => temp(17289 DOWNTO 17280) := ADC(11 DOWNTO 2);
			WHEN 1729 => temp(17299 DOWNTO 17290) := ADC(11 DOWNTO 2);
			WHEN 1730 => temp(17309 DOWNTO 17300) := ADC(11 DOWNTO 2);
			WHEN 1731 => temp(17319 DOWNTO 17310) := ADC(11 DOWNTO 2);
			WHEN 1732 => temp(17329 DOWNTO 17320) := ADC(11 DOWNTO 2);
			WHEN 1733 => temp(17339 DOWNTO 17330) := ADC(11 DOWNTO 2);
			WHEN 1734 => temp(17349 DOWNTO 17340) := ADC(11 DOWNTO 2);
			WHEN 1735 => temp(17359 DOWNTO 17350) := ADC(11 DOWNTO 2);
			WHEN 1736 => temp(17369 DOWNTO 17360) := ADC(11 DOWNTO 2);
			WHEN 1737 => temp(17379 DOWNTO 17370) := ADC(11 DOWNTO 2);
			WHEN 1738 => temp(17389 DOWNTO 17380) := ADC(11 DOWNTO 2);
			WHEN 1739 => temp(17399 DOWNTO 17390) := ADC(11 DOWNTO 2);
			WHEN 1740 => temp(17409 DOWNTO 17400) := ADC(11 DOWNTO 2);
			WHEN 1741 => temp(17419 DOWNTO 17410) := ADC(11 DOWNTO 2);
			WHEN 1742 => temp(17429 DOWNTO 17420) := ADC(11 DOWNTO 2);
			WHEN 1743 => temp(17439 DOWNTO 17430) := ADC(11 DOWNTO 2);
			WHEN 1744 => temp(17449 DOWNTO 17440) := ADC(11 DOWNTO 2);
			WHEN 1745 => temp(17459 DOWNTO 17450) := ADC(11 DOWNTO 2);
			WHEN 1746 => temp(17469 DOWNTO 17460) := ADC(11 DOWNTO 2);
			WHEN 1747 => temp(17479 DOWNTO 17470) := ADC(11 DOWNTO 2);
			WHEN 1748 => temp(17489 DOWNTO 17480) := ADC(11 DOWNTO 2);
			WHEN 1749 => temp(17499 DOWNTO 17490) := ADC(11 DOWNTO 2);
			WHEN 1750 => temp(17509 DOWNTO 17500) := ADC(11 DOWNTO 2);
			WHEN 1751 => temp(17519 DOWNTO 17510) := ADC(11 DOWNTO 2);
			WHEN 1752 => temp(17529 DOWNTO 17520) := ADC(11 DOWNTO 2);
			WHEN 1753 => temp(17539 DOWNTO 17530) := ADC(11 DOWNTO 2);
			WHEN 1754 => temp(17549 DOWNTO 17540) := ADC(11 DOWNTO 2);
			WHEN 1755 => temp(17559 DOWNTO 17550) := ADC(11 DOWNTO 2);
			WHEN 1756 => temp(17569 DOWNTO 17560) := ADC(11 DOWNTO 2);
			WHEN 1757 => temp(17579 DOWNTO 17570) := ADC(11 DOWNTO 2);
			WHEN 1758 => temp(17589 DOWNTO 17580) := ADC(11 DOWNTO 2);
			WHEN 1759 => temp(17599 DOWNTO 17590) := ADC(11 DOWNTO 2);
			WHEN 1760 => temp(17609 DOWNTO 17600) := ADC(11 DOWNTO 2);
			WHEN 1761 => temp(17619 DOWNTO 17610) := ADC(11 DOWNTO 2);
			WHEN 1762 => temp(17629 DOWNTO 17620) := ADC(11 DOWNTO 2);
			WHEN 1763 => temp(17639 DOWNTO 17630) := ADC(11 DOWNTO 2);
			WHEN 1764 => temp(17649 DOWNTO 17640) := ADC(11 DOWNTO 2);
			WHEN 1765 => temp(17659 DOWNTO 17650) := ADC(11 DOWNTO 2);
			WHEN 1766 => temp(17669 DOWNTO 17660) := ADC(11 DOWNTO 2);
			WHEN 1767 => temp(17679 DOWNTO 17670) := ADC(11 DOWNTO 2);
			WHEN 1768 => temp(17689 DOWNTO 17680) := ADC(11 DOWNTO 2);
			WHEN 1769 => temp(17699 DOWNTO 17690) := ADC(11 DOWNTO 2);
			WHEN 1770 => temp(17709 DOWNTO 17700) := ADC(11 DOWNTO 2);
			WHEN 1771 => temp(17719 DOWNTO 17710) := ADC(11 DOWNTO 2);
			WHEN 1772 => temp(17729 DOWNTO 17720) := ADC(11 DOWNTO 2);
			WHEN 1773 => temp(17739 DOWNTO 17730) := ADC(11 DOWNTO 2);
			WHEN 1774 => temp(17749 DOWNTO 17740) := ADC(11 DOWNTO 2);
			WHEN 1775 => temp(17759 DOWNTO 17750) := ADC(11 DOWNTO 2);
			WHEN 1776 => temp(17769 DOWNTO 17760) := ADC(11 DOWNTO 2);
			WHEN 1777 => temp(17779 DOWNTO 17770) := ADC(11 DOWNTO 2);
			WHEN 1778 => temp(17789 DOWNTO 17780) := ADC(11 DOWNTO 2);
			WHEN 1779 => temp(17799 DOWNTO 17790) := ADC(11 DOWNTO 2);
			WHEN 1780 => temp(17809 DOWNTO 17800) := ADC(11 DOWNTO 2);
			WHEN 1781 => temp(17819 DOWNTO 17810) := ADC(11 DOWNTO 2);
			WHEN 1782 => temp(17829 DOWNTO 17820) := ADC(11 DOWNTO 2);
			WHEN 1783 => temp(17839 DOWNTO 17830) := ADC(11 DOWNTO 2);
			WHEN 1784 => temp(17849 DOWNTO 17840) := ADC(11 DOWNTO 2);
			WHEN 1785 => temp(17859 DOWNTO 17850) := ADC(11 DOWNTO 2);
			WHEN 1786 => temp(17869 DOWNTO 17860) := ADC(11 DOWNTO 2);
			WHEN 1787 => temp(17879 DOWNTO 17870) := ADC(11 DOWNTO 2);
			WHEN 1788 => temp(17889 DOWNTO 17880) := ADC(11 DOWNTO 2);
			WHEN 1789 => temp(17899 DOWNTO 17890) := ADC(11 DOWNTO 2);
			WHEN 1790 => temp(17909 DOWNTO 17900) := ADC(11 DOWNTO 2);
			WHEN 1791 => temp(17919 DOWNTO 17910) := ADC(11 DOWNTO 2);
			WHEN 1792 => temp(17929 DOWNTO 17920) := ADC(11 DOWNTO 2);
			WHEN 1793 => temp(17939 DOWNTO 17930) := ADC(11 DOWNTO 2);
			WHEN 1794 => temp(17949 DOWNTO 17940) := ADC(11 DOWNTO 2);
			WHEN 1795 => temp(17959 DOWNTO 17950) := ADC(11 DOWNTO 2);
			WHEN 1796 => temp(17969 DOWNTO 17960) := ADC(11 DOWNTO 2);
			WHEN 1797 => temp(17979 DOWNTO 17970) := ADC(11 DOWNTO 2);
			WHEN 1798 => temp(17989 DOWNTO 17980) := ADC(11 DOWNTO 2);
			WHEN 1799 => temp(17999 DOWNTO 17990) := ADC(11 DOWNTO 2);
			WHEN 1800 => temp(18009 DOWNTO 18000) := ADC(11 DOWNTO 2);
			WHEN 1801 => temp(18019 DOWNTO 18010) := ADC(11 DOWNTO 2);
			WHEN 1802 => temp(18029 DOWNTO 18020) := ADC(11 DOWNTO 2);
			WHEN 1803 => temp(18039 DOWNTO 18030) := ADC(11 DOWNTO 2);
			WHEN 1804 => temp(18049 DOWNTO 18040) := ADC(11 DOWNTO 2);
			WHEN 1805 => temp(18059 DOWNTO 18050) := ADC(11 DOWNTO 2);
			WHEN 1806 => temp(18069 DOWNTO 18060) := ADC(11 DOWNTO 2);
			WHEN 1807 => temp(18079 DOWNTO 18070) := ADC(11 DOWNTO 2);
			WHEN 1808 => temp(18089 DOWNTO 18080) := ADC(11 DOWNTO 2);
			WHEN 1809 => temp(18099 DOWNTO 18090) := ADC(11 DOWNTO 2);
			WHEN 1810 => temp(18109 DOWNTO 18100) := ADC(11 DOWNTO 2);
			WHEN 1811 => temp(18119 DOWNTO 18110) := ADC(11 DOWNTO 2);
			WHEN 1812 => temp(18129 DOWNTO 18120) := ADC(11 DOWNTO 2);
			WHEN 1813 => temp(18139 DOWNTO 18130) := ADC(11 DOWNTO 2);
			WHEN 1814 => temp(18149 DOWNTO 18140) := ADC(11 DOWNTO 2);
			WHEN 1815 => temp(18159 DOWNTO 18150) := ADC(11 DOWNTO 2);
			WHEN 1816 => temp(18169 DOWNTO 18160) := ADC(11 DOWNTO 2);
			WHEN 1817 => temp(18179 DOWNTO 18170) := ADC(11 DOWNTO 2);
			WHEN 1818 => temp(18189 DOWNTO 18180) := ADC(11 DOWNTO 2);
			WHEN 1819 => temp(18199 DOWNTO 18190) := ADC(11 DOWNTO 2);
			WHEN 1820 => temp(18209 DOWNTO 18200) := ADC(11 DOWNTO 2);
			WHEN 1821 => temp(18219 DOWNTO 18210) := ADC(11 DOWNTO 2);
			WHEN 1822 => temp(18229 DOWNTO 18220) := ADC(11 DOWNTO 2);
			WHEN 1823 => temp(18239 DOWNTO 18230) := ADC(11 DOWNTO 2);
			WHEN 1824 => temp(18249 DOWNTO 18240) := ADC(11 DOWNTO 2);
			WHEN 1825 => temp(18259 DOWNTO 18250) := ADC(11 DOWNTO 2);
			WHEN 1826 => temp(18269 DOWNTO 18260) := ADC(11 DOWNTO 2);
			WHEN 1827 => temp(18279 DOWNTO 18270) := ADC(11 DOWNTO 2);
			WHEN 1828 => temp(18289 DOWNTO 18280) := ADC(11 DOWNTO 2);
			WHEN 1829 => temp(18299 DOWNTO 18290) := ADC(11 DOWNTO 2);
			WHEN 1830 => temp(18309 DOWNTO 18300) := ADC(11 DOWNTO 2);
			WHEN 1831 => temp(18319 DOWNTO 18310) := ADC(11 DOWNTO 2);
			WHEN 1832 => temp(18329 DOWNTO 18320) := ADC(11 DOWNTO 2);
			WHEN 1833 => temp(18339 DOWNTO 18330) := ADC(11 DOWNTO 2);
			WHEN 1834 => temp(18349 DOWNTO 18340) := ADC(11 DOWNTO 2);
			WHEN 1835 => temp(18359 DOWNTO 18350) := ADC(11 DOWNTO 2);
			WHEN 1836 => temp(18369 DOWNTO 18360) := ADC(11 DOWNTO 2);
			WHEN 1837 => temp(18379 DOWNTO 18370) := ADC(11 DOWNTO 2);
			WHEN 1838 => temp(18389 DOWNTO 18380) := ADC(11 DOWNTO 2);
			WHEN 1839 => temp(18399 DOWNTO 18390) := ADC(11 DOWNTO 2);
			WHEN 1840 => temp(18409 DOWNTO 18400) := ADC(11 DOWNTO 2);
			WHEN 1841 => temp(18419 DOWNTO 18410) := ADC(11 DOWNTO 2);
			WHEN 1842 => temp(18429 DOWNTO 18420) := ADC(11 DOWNTO 2);
			WHEN 1843 => temp(18439 DOWNTO 18430) := ADC(11 DOWNTO 2);
			WHEN 1844 => temp(18449 DOWNTO 18440) := ADC(11 DOWNTO 2);
			WHEN 1845 => temp(18459 DOWNTO 18450) := ADC(11 DOWNTO 2);
			WHEN 1846 => temp(18469 DOWNTO 18460) := ADC(11 DOWNTO 2);
			WHEN 1847 => temp(18479 DOWNTO 18470) := ADC(11 DOWNTO 2);
			WHEN 1848 => temp(18489 DOWNTO 18480) := ADC(11 DOWNTO 2);
			WHEN 1849 => temp(18499 DOWNTO 18490) := ADC(11 DOWNTO 2);
			WHEN 1850 => temp(18509 DOWNTO 18500) := ADC(11 DOWNTO 2);
			WHEN 1851 => temp(18519 DOWNTO 18510) := ADC(11 DOWNTO 2);
			WHEN 1852 => temp(18529 DOWNTO 18520) := ADC(11 DOWNTO 2);
			WHEN 1853 => temp(18539 DOWNTO 18530) := ADC(11 DOWNTO 2);
			WHEN 1854 => temp(18549 DOWNTO 18540) := ADC(11 DOWNTO 2);
			WHEN 1855 => temp(18559 DOWNTO 18550) := ADC(11 DOWNTO 2);
			WHEN 1856 => temp(18569 DOWNTO 18560) := ADC(11 DOWNTO 2);
			WHEN 1857 => temp(18579 DOWNTO 18570) := ADC(11 DOWNTO 2);
			WHEN 1858 => temp(18589 DOWNTO 18580) := ADC(11 DOWNTO 2);
			WHEN 1859 => temp(18599 DOWNTO 18590) := ADC(11 DOWNTO 2);
			WHEN 1860 => temp(18609 DOWNTO 18600) := ADC(11 DOWNTO 2);
			WHEN 1861 => temp(18619 DOWNTO 18610) := ADC(11 DOWNTO 2);
			WHEN 1862 => temp(18629 DOWNTO 18620) := ADC(11 DOWNTO 2);
			WHEN 1863 => temp(18639 DOWNTO 18630) := ADC(11 DOWNTO 2);
			WHEN 1864 => temp(18649 DOWNTO 18640) := ADC(11 DOWNTO 2);
			WHEN 1865 => temp(18659 DOWNTO 18650) := ADC(11 DOWNTO 2);
			WHEN 1866 => temp(18669 DOWNTO 18660) := ADC(11 DOWNTO 2);
			WHEN 1867 => temp(18679 DOWNTO 18670) := ADC(11 DOWNTO 2);
			WHEN 1868 => temp(18689 DOWNTO 18680) := ADC(11 DOWNTO 2);
			WHEN 1869 => temp(18699 DOWNTO 18690) := ADC(11 DOWNTO 2);
			WHEN 1870 => temp(18709 DOWNTO 18700) := ADC(11 DOWNTO 2);
			WHEN 1871 => temp(18719 DOWNTO 18710) := ADC(11 DOWNTO 2);
			WHEN 1872 => temp(18729 DOWNTO 18720) := ADC(11 DOWNTO 2);
			WHEN 1873 => temp(18739 DOWNTO 18730) := ADC(11 DOWNTO 2);
			WHEN 1874 => temp(18749 DOWNTO 18740) := ADC(11 DOWNTO 2);
			WHEN 1875 => temp(18759 DOWNTO 18750) := ADC(11 DOWNTO 2);
			WHEN 1876 => temp(18769 DOWNTO 18760) := ADC(11 DOWNTO 2);
			WHEN 1877 => temp(18779 DOWNTO 18770) := ADC(11 DOWNTO 2);
			WHEN 1878 => temp(18789 DOWNTO 18780) := ADC(11 DOWNTO 2);
			WHEN 1879 => temp(18799 DOWNTO 18790) := ADC(11 DOWNTO 2);
			WHEN 1880 => temp(18809 DOWNTO 18800) := ADC(11 DOWNTO 2);
			WHEN 1881 => temp(18819 DOWNTO 18810) := ADC(11 DOWNTO 2);
			WHEN 1882 => temp(18829 DOWNTO 18820) := ADC(11 DOWNTO 2);
			WHEN 1883 => temp(18839 DOWNTO 18830) := ADC(11 DOWNTO 2);
			WHEN 1884 => temp(18849 DOWNTO 18840) := ADC(11 DOWNTO 2);
			WHEN 1885 => temp(18859 DOWNTO 18850) := ADC(11 DOWNTO 2);
			WHEN 1886 => temp(18869 DOWNTO 18860) := ADC(11 DOWNTO 2);
			WHEN 1887 => temp(18879 DOWNTO 18870) := ADC(11 DOWNTO 2);
			WHEN 1888 => temp(18889 DOWNTO 18880) := ADC(11 DOWNTO 2);
			WHEN 1889 => temp(18899 DOWNTO 18890) := ADC(11 DOWNTO 2);
			WHEN 1890 => temp(18909 DOWNTO 18900) := ADC(11 DOWNTO 2);
			WHEN 1891 => temp(18919 DOWNTO 18910) := ADC(11 DOWNTO 2);
			WHEN 1892 => temp(18929 DOWNTO 18920) := ADC(11 DOWNTO 2);
			WHEN 1893 => temp(18939 DOWNTO 18930) := ADC(11 DOWNTO 2);
			WHEN 1894 => temp(18949 DOWNTO 18940) := ADC(11 DOWNTO 2);
			WHEN 1895 => temp(18959 DOWNTO 18950) := ADC(11 DOWNTO 2);
			WHEN 1896 => temp(18969 DOWNTO 18960) := ADC(11 DOWNTO 2);
			WHEN 1897 => temp(18979 DOWNTO 18970) := ADC(11 DOWNTO 2);
			WHEN 1898 => temp(18989 DOWNTO 18980) := ADC(11 DOWNTO 2);
			WHEN 1899 => temp(18999 DOWNTO 18990) := ADC(11 DOWNTO 2);
			WHEN 1900 => temp(19009 DOWNTO 19000) := ADC(11 DOWNTO 2);
			WHEN 1901 => temp(19019 DOWNTO 19010) := ADC(11 DOWNTO 2);
			WHEN 1902 => temp(19029 DOWNTO 19020) := ADC(11 DOWNTO 2);
			WHEN 1903 => temp(19039 DOWNTO 19030) := ADC(11 DOWNTO 2);
			WHEN 1904 => temp(19049 DOWNTO 19040) := ADC(11 DOWNTO 2);
			WHEN 1905 => temp(19059 DOWNTO 19050) := ADC(11 DOWNTO 2);
			WHEN 1906 => temp(19069 DOWNTO 19060) := ADC(11 DOWNTO 2);
			WHEN 1907 => temp(19079 DOWNTO 19070) := ADC(11 DOWNTO 2);
			WHEN 1908 => temp(19089 DOWNTO 19080) := ADC(11 DOWNTO 2);
			WHEN 1909 => temp(19099 DOWNTO 19090) := ADC(11 DOWNTO 2);
			WHEN 1910 => temp(19109 DOWNTO 19100) := ADC(11 DOWNTO 2);
			WHEN 1911 => temp(19119 DOWNTO 19110) := ADC(11 DOWNTO 2);
			WHEN 1912 => temp(19129 DOWNTO 19120) := ADC(11 DOWNTO 2);
			WHEN 1913 => temp(19139 DOWNTO 19130) := ADC(11 DOWNTO 2);
			WHEN 1914 => temp(19149 DOWNTO 19140) := ADC(11 DOWNTO 2);
			WHEN 1915 => temp(19159 DOWNTO 19150) := ADC(11 DOWNTO 2);
			WHEN 1916 => temp(19169 DOWNTO 19160) := ADC(11 DOWNTO 2);
			WHEN 1917 => temp(19179 DOWNTO 19170) := ADC(11 DOWNTO 2);
			WHEN 1918 => temp(19189 DOWNTO 19180) := ADC(11 DOWNTO 2);
			WHEN 1919 => temp(19199 DOWNTO 19190) := ADC(11 DOWNTO 2);
			WHEN 1920 => temp(19209 DOWNTO 19200) := ADC(11 DOWNTO 2);
			WHEN 1921 => temp(19219 DOWNTO 19210) := ADC(11 DOWNTO 2);
			WHEN 1922 => temp(19229 DOWNTO 19220) := ADC(11 DOWNTO 2);
			WHEN 1923 => temp(19239 DOWNTO 19230) := ADC(11 DOWNTO 2);
			WHEN 1924 => temp(19249 DOWNTO 19240) := ADC(11 DOWNTO 2);
			WHEN 1925 => temp(19259 DOWNTO 19250) := ADC(11 DOWNTO 2);
			WHEN 1926 => temp(19269 DOWNTO 19260) := ADC(11 DOWNTO 2);
			WHEN 1927 => temp(19279 DOWNTO 19270) := ADC(11 DOWNTO 2);
			WHEN 1928 => temp(19289 DOWNTO 19280) := ADC(11 DOWNTO 2);
			WHEN 1929 => temp(19299 DOWNTO 19290) := ADC(11 DOWNTO 2);
			WHEN 1930 => temp(19309 DOWNTO 19300) := ADC(11 DOWNTO 2);
			WHEN 1931 => temp(19319 DOWNTO 19310) := ADC(11 DOWNTO 2);
			WHEN 1932 => temp(19329 DOWNTO 19320) := ADC(11 DOWNTO 2);
			WHEN 1933 => temp(19339 DOWNTO 19330) := ADC(11 DOWNTO 2);
			WHEN 1934 => temp(19349 DOWNTO 19340) := ADC(11 DOWNTO 2);
			WHEN 1935 => temp(19359 DOWNTO 19350) := ADC(11 DOWNTO 2);
			WHEN 1936 => temp(19369 DOWNTO 19360) := ADC(11 DOWNTO 2);
			WHEN 1937 => temp(19379 DOWNTO 19370) := ADC(11 DOWNTO 2);
			WHEN 1938 => temp(19389 DOWNTO 19380) := ADC(11 DOWNTO 2);
			WHEN 1939 => temp(19399 DOWNTO 19390) := ADC(11 DOWNTO 2);
			WHEN 1940 => temp(19409 DOWNTO 19400) := ADC(11 DOWNTO 2);
			WHEN 1941 => temp(19419 DOWNTO 19410) := ADC(11 DOWNTO 2);
			WHEN 1942 => temp(19429 DOWNTO 19420) := ADC(11 DOWNTO 2);
			WHEN 1943 => temp(19439 DOWNTO 19430) := ADC(11 DOWNTO 2);
			WHEN 1944 => temp(19449 DOWNTO 19440) := ADC(11 DOWNTO 2);
			WHEN 1945 => temp(19459 DOWNTO 19450) := ADC(11 DOWNTO 2);
			WHEN 1946 => temp(19469 DOWNTO 19460) := ADC(11 DOWNTO 2);
			WHEN 1947 => temp(19479 DOWNTO 19470) := ADC(11 DOWNTO 2);
			WHEN 1948 => temp(19489 DOWNTO 19480) := ADC(11 DOWNTO 2);
			WHEN 1949 => temp(19499 DOWNTO 19490) := ADC(11 DOWNTO 2);
			WHEN 1950 => temp(19509 DOWNTO 19500) := ADC(11 DOWNTO 2);
			WHEN 1951 => temp(19519 DOWNTO 19510) := ADC(11 DOWNTO 2);
			WHEN 1952 => temp(19529 DOWNTO 19520) := ADC(11 DOWNTO 2);
			WHEN 1953 => temp(19539 DOWNTO 19530) := ADC(11 DOWNTO 2);
			WHEN 1954 => temp(19549 DOWNTO 19540) := ADC(11 DOWNTO 2);
			WHEN 1955 => temp(19559 DOWNTO 19550) := ADC(11 DOWNTO 2);
			WHEN 1956 => temp(19569 DOWNTO 19560) := ADC(11 DOWNTO 2);
			WHEN 1957 => temp(19579 DOWNTO 19570) := ADC(11 DOWNTO 2);
			WHEN 1958 => temp(19589 DOWNTO 19580) := ADC(11 DOWNTO 2);
			WHEN 1959 => temp(19599 DOWNTO 19590) := ADC(11 DOWNTO 2);
			WHEN 1960 => temp(19609 DOWNTO 19600) := ADC(11 DOWNTO 2);
			WHEN 1961 => temp(19619 DOWNTO 19610) := ADC(11 DOWNTO 2);
			WHEN 1962 => temp(19629 DOWNTO 19620) := ADC(11 DOWNTO 2);
			WHEN 1963 => temp(19639 DOWNTO 19630) := ADC(11 DOWNTO 2);
			WHEN 1964 => temp(19649 DOWNTO 19640) := ADC(11 DOWNTO 2);
			WHEN 1965 => temp(19659 DOWNTO 19650) := ADC(11 DOWNTO 2);
			WHEN 1966 => temp(19669 DOWNTO 19660) := ADC(11 DOWNTO 2);
			WHEN 1967 => temp(19679 DOWNTO 19670) := ADC(11 DOWNTO 2);
			WHEN 1968 => temp(19689 DOWNTO 19680) := ADC(11 DOWNTO 2);
			WHEN 1969 => temp(19699 DOWNTO 19690) := ADC(11 DOWNTO 2);
			WHEN 1970 => temp(19709 DOWNTO 19700) := ADC(11 DOWNTO 2);
			WHEN 1971 => temp(19719 DOWNTO 19710) := ADC(11 DOWNTO 2);
			WHEN 1972 => temp(19729 DOWNTO 19720) := ADC(11 DOWNTO 2);
			WHEN 1973 => temp(19739 DOWNTO 19730) := ADC(11 DOWNTO 2);
			WHEN 1974 => temp(19749 DOWNTO 19740) := ADC(11 DOWNTO 2);
			WHEN 1975 => temp(19759 DOWNTO 19750) := ADC(11 DOWNTO 2);
			WHEN 1976 => temp(19769 DOWNTO 19760) := ADC(11 DOWNTO 2);
			WHEN 1977 => temp(19779 DOWNTO 19770) := ADC(11 DOWNTO 2);
			WHEN 1978 => temp(19789 DOWNTO 19780) := ADC(11 DOWNTO 2);
			WHEN 1979 => temp(19799 DOWNTO 19790) := ADC(11 DOWNTO 2);
			WHEN 1980 => temp(19809 DOWNTO 19800) := ADC(11 DOWNTO 2);
			WHEN 1981 => temp(19819 DOWNTO 19810) := ADC(11 DOWNTO 2);
			WHEN 1982 => temp(19829 DOWNTO 19820) := ADC(11 DOWNTO 2);
			WHEN 1983 => temp(19839 DOWNTO 19830) := ADC(11 DOWNTO 2);
			WHEN 1984 => temp(19849 DOWNTO 19840) := ADC(11 DOWNTO 2);
			WHEN 1985 => temp(19859 DOWNTO 19850) := ADC(11 DOWNTO 2);
			WHEN 1986 => temp(19869 DOWNTO 19860) := ADC(11 DOWNTO 2);
			WHEN 1987 => temp(19879 DOWNTO 19870) := ADC(11 DOWNTO 2);
			WHEN 1988 => temp(19889 DOWNTO 19880) := ADC(11 DOWNTO 2);
			WHEN 1989 => temp(19899 DOWNTO 19890) := ADC(11 DOWNTO 2);
			WHEN 1990 => temp(19909 DOWNTO 19900) := ADC(11 DOWNTO 2);
			WHEN 1991 => temp(19919 DOWNTO 19910) := ADC(11 DOWNTO 2);
			WHEN 1992 => temp(19929 DOWNTO 19920) := ADC(11 DOWNTO 2);
			WHEN 1993 => temp(19939 DOWNTO 19930) := ADC(11 DOWNTO 2);
			WHEN 1994 => temp(19949 DOWNTO 19940) := ADC(11 DOWNTO 2);
			WHEN 1995 => temp(19959 DOWNTO 19950) := ADC(11 DOWNTO 2);
			WHEN 1996 => temp(19969 DOWNTO 19960) := ADC(11 DOWNTO 2);
			WHEN 1997 => temp(19979 DOWNTO 19970) := ADC(11 DOWNTO 2);
			WHEN 1998 => temp(19989 DOWNTO 19980) := ADC(11 DOWNTO 2);
			WHEN 1999 => temp(19999 DOWNTO 19990) := ADC(11 DOWNTO 2);
			WHEN 2000 => temp(20009 DOWNTO 20000) := ADC(11 DOWNTO 2);
			WHEN 2001 => temp(20019 DOWNTO 20010) := ADC(11 DOWNTO 2);
			WHEN 2002 => temp(20029 DOWNTO 20020) := ADC(11 DOWNTO 2);
			WHEN 2003 => temp(20039 DOWNTO 20030) := ADC(11 DOWNTO 2);
			WHEN 2004 => temp(20049 DOWNTO 20040) := ADC(11 DOWNTO 2);
			WHEN 2005 => temp(20059 DOWNTO 20050) := ADC(11 DOWNTO 2);
			WHEN 2006 => temp(20069 DOWNTO 20060) := ADC(11 DOWNTO 2);
			WHEN 2007 => temp(20079 DOWNTO 20070) := ADC(11 DOWNTO 2);
			WHEN 2008 => temp(20089 DOWNTO 20080) := ADC(11 DOWNTO 2);
			WHEN 2009 => temp(20099 DOWNTO 20090) := ADC(11 DOWNTO 2);
			WHEN 2010 => temp(20109 DOWNTO 20100) := ADC(11 DOWNTO 2);
			WHEN 2011 => temp(20119 DOWNTO 20110) := ADC(11 DOWNTO 2);
			WHEN 2012 => temp(20129 DOWNTO 20120) := ADC(11 DOWNTO 2);
			WHEN 2013 => temp(20139 DOWNTO 20130) := ADC(11 DOWNTO 2);
			WHEN 2014 => temp(20149 DOWNTO 20140) := ADC(11 DOWNTO 2);
			WHEN 2015 => temp(20159 DOWNTO 20150) := ADC(11 DOWNTO 2);
			WHEN 2016 => temp(20169 DOWNTO 20160) := ADC(11 DOWNTO 2);
			WHEN 2017 => temp(20179 DOWNTO 20170) := ADC(11 DOWNTO 2);
			WHEN 2018 => temp(20189 DOWNTO 20180) := ADC(11 DOWNTO 2);
			WHEN 2019 => temp(20199 DOWNTO 20190) := ADC(11 DOWNTO 2);
			WHEN 2020 => temp(20209 DOWNTO 20200) := ADC(11 DOWNTO 2);
			WHEN 2021 => temp(20219 DOWNTO 20210) := ADC(11 DOWNTO 2);
			WHEN 2022 => temp(20229 DOWNTO 20220) := ADC(11 DOWNTO 2);
			WHEN 2023 => temp(20239 DOWNTO 20230) := ADC(11 DOWNTO 2);
			WHEN 2024 => temp(20249 DOWNTO 20240) := ADC(11 DOWNTO 2);
			WHEN 2025 => temp(20259 DOWNTO 20250) := ADC(11 DOWNTO 2);
			WHEN 2026 => temp(20269 DOWNTO 20260) := ADC(11 DOWNTO 2);
			WHEN 2027 => temp(20279 DOWNTO 20270) := ADC(11 DOWNTO 2);
			WHEN 2028 => temp(20289 DOWNTO 20280) := ADC(11 DOWNTO 2);
			WHEN 2029 => temp(20299 DOWNTO 20290) := ADC(11 DOWNTO 2);
			WHEN 2030 => temp(20309 DOWNTO 20300) := ADC(11 DOWNTO 2);
			WHEN 2031 => temp(20319 DOWNTO 20310) := ADC(11 DOWNTO 2);
			WHEN 2032 => temp(20329 DOWNTO 20320) := ADC(11 DOWNTO 2);
			WHEN 2033 => temp(20339 DOWNTO 20330) := ADC(11 DOWNTO 2);
			WHEN 2034 => temp(20349 DOWNTO 20340) := ADC(11 DOWNTO 2);
			WHEN 2035 => temp(20359 DOWNTO 20350) := ADC(11 DOWNTO 2);
			WHEN 2036 => temp(20369 DOWNTO 20360) := ADC(11 DOWNTO 2);
			WHEN 2037 => temp(20379 DOWNTO 20370) := ADC(11 DOWNTO 2);
			WHEN 2038 => temp(20389 DOWNTO 20380) := ADC(11 DOWNTO 2);
			WHEN 2039 => temp(20399 DOWNTO 20390) := ADC(11 DOWNTO 2);
			WHEN 2040 => temp(20409 DOWNTO 20400) := ADC(11 DOWNTO 2);
			WHEN 2041 => temp(20419 DOWNTO 20410) := ADC(11 DOWNTO 2);
			WHEN 2042 => temp(20429 DOWNTO 20420) := ADC(11 DOWNTO 2);
			WHEN 2043 => temp(20439 DOWNTO 20430) := ADC(11 DOWNTO 2);
			WHEN 2044 => temp(20449 DOWNTO 20440) := ADC(11 DOWNTO 2);
			WHEN 2045 => temp(20459 DOWNTO 20450) := ADC(11 DOWNTO 2);
			WHEN 2046 => temp(20469 DOWNTO 20460) := ADC(11 DOWNTO 2);
			WHEN 2047 => temp(20479 DOWNTO 20470) := ADC(11 DOWNTO 2);		
			WHEN OTHERS => NULL;
				END CASE;
			done <= '1';
		ELSE 
			done <= '0';
		END IF;
		samples <= temp;
	END IF;
	END PROCESS;
END;