// nios2VGA.v

// Generated using ACDS version 13.0sp1 232 at 2014.02.02.13:03:56

`timescale 1 ps / 1 ps
module nios2VGA (
		input  wire        clk_clk,                                  //                               clk.clk
		input  wire        reset_reset_n,                            //                             reset.reset_n
		output wire [17:0] red_led_pio_external_connection_export,   //   red_led_pio_external_connection.export
		output wire        vga_controller_external_CLK,              //           vga_controller_external.CLK
		output wire        vga_controller_external_HS,               //                                  .HS
		output wire        vga_controller_external_VS,               //                                  .VS
		output wire        vga_controller_external_BLANK,            //                                  .BLANK
		output wire        vga_controller_external_SYNC,             //                                  .SYNC
		output wire [9:0]  vga_controller_external_R,                //                                  .R
		output wire [9:0]  vga_controller_external_G,                //                                  .G
		output wire [9:0]  vga_controller_external_B,                //                                  .B
		inout  wire [15:0] sram_external_interface_DQ,               //           sram_external_interface.DQ
		output wire [17:0] sram_external_interface_ADDR,             //                                  .ADDR
		output wire        sram_external_interface_LB_N,             //                                  .LB_N
		output wire        sram_external_interface_UB_N,             //                                  .UB_N
		output wire        sram_external_interface_CE_N,             //                                  .CE_N
		output wire        sram_external_interface_OE_N,             //                                  .OE_N
		output wire        sram_external_interface_WE_N,             //                                  .WE_N
		output wire        vga_clock_out_clk_clk,                    //                 vga_clock_out_clk.clk
		output wire [8:0]  green_led_pio_external_connection_export, // green_led_pio_external_connection.export
		output wire        sdram_clock_clk,                          //                       sdram_clock.clk
		input  wire [7:0]  nios_cntrl_in_export,                     //                     nios_cntrl_in.export
		output wire [7:0]  nios_cntrl_out_export,                    //                    nios_cntrl_out.export
		input  wire [31:0] fft_in_0_export,                          //                          fft_in_0.export
		input  wire [31:0] fft_in_1_export,                          //                          fft_in_1.export
		input  wire [31:0] fft_in_2_export,                          //                          fft_in_2.export
		input  wire [31:0] fft_in_3_export,                          //                          fft_in_3.export
		input  wire [7:0]  rotary_in_export,                         //                         rotary_in.export
		input  wire [31:0] fft_in_4_export,                          //                          fft_in_4.export
		input  wire [31:0] fft_in_5_export,                          //                          fft_in_5.export
		input  wire [31:0] fft_in_6_export,                          //                          fft_in_6.export
		input  wire [31:0] fft_in_7_export                           //                          fft_in_7.export
	);

	wire          external_clocks_sys_clk_clk;                                                                                         // external_clocks:sys_clk -> [Alpha_Blending:clk, SRAM:clk, SRAM_avalon_sram_slave_translator:clk, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Character_buffer:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Character_buffer_avalon_char_control_slave_translator:clk, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:clk, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Dual_Clock_FIFO:clk_stream_in, VGA_Pixel_Buffer:clk, VGA_Pixel_Buffer_avalon_control_slave_translator:clk, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:clk, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, VGA_Scaler:clk, VGA_pixel_RGB_Resampler:clk, addr_router_001:clk, burst_adapter:clk, burst_adapter_001:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux_001:clk, crosser:out_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, crosser_004:out_clk, crosser_005:out_clk, crosser_006:out_clk, crosser_007:in_clk, crosser_008:in_clk, crosser_009:in_clk, id_router_001:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rst_controller_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk]
	wire          vga_character_buffer_avalon_char_source_endofpacket;                                                                 // VGA_Character_buffer:stream_endofpacket -> Alpha_Blending:foreground_endofpacket
	wire          vga_character_buffer_avalon_char_source_valid;                                                                       // VGA_Character_buffer:stream_valid -> Alpha_Blending:foreground_valid
	wire          vga_character_buffer_avalon_char_source_startofpacket;                                                               // VGA_Character_buffer:stream_startofpacket -> Alpha_Blending:foreground_startofpacket
	wire   [39:0] vga_character_buffer_avalon_char_source_data;                                                                        // VGA_Character_buffer:stream_data -> Alpha_Blending:foreground_data
	wire          vga_character_buffer_avalon_char_source_ready;                                                                       // Alpha_Blending:foreground_ready -> VGA_Character_buffer:stream_ready
	wire          alpha_blending_avalon_blended_source_endofpacket;                                                                    // Alpha_Blending:output_endofpacket -> VGA_Dual_Clock_FIFO:stream_in_endofpacket
	wire          alpha_blending_avalon_blended_source_valid;                                                                          // Alpha_Blending:output_valid -> VGA_Dual_Clock_FIFO:stream_in_valid
	wire          alpha_blending_avalon_blended_source_startofpacket;                                                                  // Alpha_Blending:output_startofpacket -> VGA_Dual_Clock_FIFO:stream_in_startofpacket
	wire   [29:0] alpha_blending_avalon_blended_source_data;                                                                           // Alpha_Blending:output_data -> VGA_Dual_Clock_FIFO:stream_in_data
	wire          alpha_blending_avalon_blended_source_ready;                                                                          // VGA_Dual_Clock_FIFO:stream_in_ready -> Alpha_Blending:output_ready
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                                                             // VGA_Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_valid;                                                                   // VGA_Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                                                           // VGA_Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire   [29:0] vga_dual_clock_fifo_avalon_dc_buffer_source_data;                                                                    // VGA_Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_ready;                                                                   // VGA_Controller:ready -> VGA_Dual_Clock_FIFO:stream_out_ready
	wire          vga_scaler_avalon_scaler_source_endofpacket;                                                                         // VGA_Scaler:stream_out_endofpacket -> Alpha_Blending:background_endofpacket
	wire          vga_scaler_avalon_scaler_source_valid;                                                                               // VGA_Scaler:stream_out_valid -> Alpha_Blending:background_valid
	wire          vga_scaler_avalon_scaler_source_startofpacket;                                                                       // VGA_Scaler:stream_out_startofpacket -> Alpha_Blending:background_startofpacket
	wire   [29:0] vga_scaler_avalon_scaler_source_data;                                                                                // VGA_Scaler:stream_out_data -> Alpha_Blending:background_data
	wire          vga_scaler_avalon_scaler_source_ready;                                                                               // Alpha_Blending:background_ready -> VGA_Scaler:stream_out_ready
	wire          vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket;                                                               // VGA_pixel_RGB_Resampler:stream_out_endofpacket -> VGA_Scaler:stream_in_endofpacket
	wire          vga_pixel_rgb_resampler_avalon_rgb_source_valid;                                                                     // VGA_pixel_RGB_Resampler:stream_out_valid -> VGA_Scaler:stream_in_valid
	wire          vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket;                                                             // VGA_pixel_RGB_Resampler:stream_out_startofpacket -> VGA_Scaler:stream_in_startofpacket
	wire   [29:0] vga_pixel_rgb_resampler_avalon_rgb_source_data;                                                                      // VGA_pixel_RGB_Resampler:stream_out_data -> VGA_Scaler:stream_in_data
	wire          vga_pixel_rgb_resampler_avalon_rgb_source_ready;                                                                     // VGA_Scaler:stream_in_ready -> VGA_pixel_RGB_Resampler:stream_out_ready
	wire          vga_pixel_buffer_avalon_pixel_source_endofpacket;                                                                    // VGA_Pixel_Buffer:stream_endofpacket -> VGA_pixel_RGB_Resampler:stream_in_endofpacket
	wire          vga_pixel_buffer_avalon_pixel_source_valid;                                                                          // VGA_Pixel_Buffer:stream_valid -> VGA_pixel_RGB_Resampler:stream_in_valid
	wire          vga_pixel_buffer_avalon_pixel_source_startofpacket;                                                                  // VGA_Pixel_Buffer:stream_startofpacket -> VGA_pixel_RGB_Resampler:stream_in_startofpacket
	wire   [15:0] vga_pixel_buffer_avalon_pixel_source_data;                                                                           // VGA_Pixel_Buffer:stream_data -> VGA_pixel_RGB_Resampler:stream_in_data
	wire          vga_pixel_buffer_avalon_pixel_source_ready;                                                                          // VGA_pixel_RGB_Resampler:stream_in_ready -> VGA_Pixel_Buffer:stream_ready
	wire          cpu_instruction_master_waitrequest;                                                                                  // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [19:0] cpu_instruction_master_address;                                                                                      // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                                         // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                                     // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          vga_pixel_buffer_avalon_pixel_dma_master_waitrequest;                                                                // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_waitrequest -> VGA_Pixel_Buffer:master_waitrequest
	wire   [31:0] vga_pixel_buffer_avalon_pixel_dma_master_address;                                                                    // VGA_Pixel_Buffer:master_address -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_address
	wire          vga_pixel_buffer_avalon_pixel_dma_master_lock;                                                                       // VGA_Pixel_Buffer:master_arbiterlock -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_lock
	wire          vga_pixel_buffer_avalon_pixel_dma_master_read;                                                                       // VGA_Pixel_Buffer:master_read -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_read
	wire   [15:0] vga_pixel_buffer_avalon_pixel_dma_master_readdata;                                                                   // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_readdata -> VGA_Pixel_Buffer:master_readdata
	wire          vga_pixel_buffer_avalon_pixel_dma_master_readdatavalid;                                                              // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:av_readdatavalid -> VGA_Pixel_Buffer:master_readdatavalid
	wire          cpu_data_master_waitrequest;                                                                                         // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                                           // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [19:0] cpu_data_master_address;                                                                                             // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                               // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                                // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                                            // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                                         // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire    [3:0] cpu_data_master_byteenable;                                                                                          // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                                    // cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                      // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                        // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                          // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                                           // cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                       // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                                    // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                     // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                                     // SRAM_avalon_sram_slave_translator:av_writedata -> SRAM:writedata
	wire   [17:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                                       // SRAM_avalon_sram_slave_translator:av_address -> SRAM:address
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                                         // SRAM_avalon_sram_slave_translator:av_write -> SRAM:write
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                                          // SRAM_avalon_sram_slave_translator:av_read -> SRAM:read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                                      // SRAM:readdata -> SRAM_avalon_sram_slave_translator:av_readdata
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                                 // SRAM:readdatavalid -> SRAM_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                                    // SRAM_avalon_sram_slave_translator:av_byteenable -> SRAM:byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                              // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                                // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                                  // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                               // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                                    // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                     // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                                 // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata;                                                           // sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	wire    [2:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_address;                                                             // sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                          // sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_write;                                                               // sys_clk_timer_s1_translator:av_write -> sys_clk_timer:write_n
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata;                                                            // sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                                          // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                                         // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] red_led_pio_s1_translator_avalon_anti_slave_0_writedata;                                                             // red_led_pio_s1_translator:av_writedata -> red_led_pio:writedata
	wire    [1:0] red_led_pio_s1_translator_avalon_anti_slave_0_address;                                                               // red_led_pio_s1_translator:av_address -> red_led_pio:address
	wire          red_led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                            // red_led_pio_s1_translator:av_chipselect -> red_led_pio:chipselect
	wire          red_led_pio_s1_translator_avalon_anti_slave_0_write;                                                                 // red_led_pio_s1_translator:av_write -> red_led_pio:write_n
	wire   [31:0] red_led_pio_s1_translator_avalon_anti_slave_0_readdata;                                                              // red_led_pio:readdata -> red_led_pio_s1_translator:av_readdata
	wire   [31:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata;                             // VGA_Character_buffer_avalon_char_control_slave_translator:av_writedata -> VGA_Character_buffer:ctrl_writedata
	wire    [0:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address;                               // VGA_Character_buffer_avalon_char_control_slave_translator:av_address -> VGA_Character_buffer:ctrl_address
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect;                            // VGA_Character_buffer_avalon_char_control_slave_translator:av_chipselect -> VGA_Character_buffer:ctrl_chipselect
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write;                                 // VGA_Character_buffer_avalon_char_control_slave_translator:av_write -> VGA_Character_buffer:ctrl_write
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read;                                  // VGA_Character_buffer_avalon_char_control_slave_translator:av_read -> VGA_Character_buffer:ctrl_read
	wire   [31:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata;                              // VGA_Character_buffer:ctrl_readdata -> VGA_Character_buffer_avalon_char_control_slave_translator:av_readdata
	wire    [3:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable;                            // VGA_Character_buffer_avalon_char_control_slave_translator:av_byteenable -> VGA_Character_buffer:ctrl_byteenable
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest;                            // VGA_Character_buffer:buf_waitrequest -> VGA_Character_buffer_avalon_char_buffer_slave_translator:av_waitrequest
	wire    [7:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata;                              // VGA_Character_buffer_avalon_char_buffer_slave_translator:av_writedata -> VGA_Character_buffer:buf_writedata
	wire   [12:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address;                                // VGA_Character_buffer_avalon_char_buffer_slave_translator:av_address -> VGA_Character_buffer:buf_address
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect;                             // VGA_Character_buffer_avalon_char_buffer_slave_translator:av_chipselect -> VGA_Character_buffer:buf_chipselect
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write;                                  // VGA_Character_buffer_avalon_char_buffer_slave_translator:av_write -> VGA_Character_buffer:buf_write
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read;                                   // VGA_Character_buffer_avalon_char_buffer_slave_translator:av_read -> VGA_Character_buffer:buf_read
	wire    [7:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata;                               // VGA_Character_buffer:buf_readdata -> VGA_Character_buffer_avalon_char_buffer_slave_translator:av_readdata
	wire    [0:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable;                             // VGA_Character_buffer_avalon_char_buffer_slave_translator:av_byteenable -> VGA_Character_buffer:buf_byteenable
	wire   [31:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_writedata;                                      // VGA_Pixel_Buffer_avalon_control_slave_translator:av_writedata -> VGA_Pixel_Buffer:slave_writedata
	wire    [1:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_address;                                        // VGA_Pixel_Buffer_avalon_control_slave_translator:av_address -> VGA_Pixel_Buffer:slave_address
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_write;                                          // VGA_Pixel_Buffer_avalon_control_slave_translator:av_write -> VGA_Pixel_Buffer:slave_write
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_read;                                           // VGA_Pixel_Buffer_avalon_control_slave_translator:av_read -> VGA_Pixel_Buffer:slave_read
	wire   [31:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_readdata;                                       // VGA_Pixel_Buffer:slave_readdata -> VGA_Pixel_Buffer_avalon_control_slave_translator:av_readdata
	wire    [3:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_byteenable;                                     // VGA_Pixel_Buffer_avalon_control_slave_translator:av_byteenable -> VGA_Pixel_Buffer:slave_byteenable
	wire   [31:0] green_led_pio_s1_translator_avalon_anti_slave_0_writedata;                                                           // green_led_pio_s1_translator:av_writedata -> green_led_pio:writedata
	wire    [1:0] green_led_pio_s1_translator_avalon_anti_slave_0_address;                                                             // green_led_pio_s1_translator:av_address -> green_led_pio:address
	wire          green_led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                          // green_led_pio_s1_translator:av_chipselect -> green_led_pio:chipselect
	wire          green_led_pio_s1_translator_avalon_anti_slave_0_write;                                                               // green_led_pio_s1_translator:av_write -> green_led_pio:write_n
	wire   [31:0] green_led_pio_s1_translator_avalon_anti_slave_0_readdata;                                                            // green_led_pio:readdata -> green_led_pio_s1_translator:av_readdata
	wire    [1:0] control_in_s1_translator_avalon_anti_slave_0_address;                                                                // control_in_s1_translator:av_address -> control_in:address
	wire   [31:0] control_in_s1_translator_avalon_anti_slave_0_readdata;                                                               // control_in:readdata -> control_in_s1_translator:av_readdata
	wire   [31:0] control_out_s1_translator_avalon_anti_slave_0_writedata;                                                             // control_out_s1_translator:av_writedata -> control_out:writedata
	wire    [1:0] control_out_s1_translator_avalon_anti_slave_0_address;                                                               // control_out_s1_translator:av_address -> control_out:address
	wire          control_out_s1_translator_avalon_anti_slave_0_chipselect;                                                            // control_out_s1_translator:av_chipselect -> control_out:chipselect
	wire          control_out_s1_translator_avalon_anti_slave_0_write;                                                                 // control_out_s1_translator:av_write -> control_out:write_n
	wire   [31:0] control_out_s1_translator_avalon_anti_slave_0_readdata;                                                              // control_out:readdata -> control_out_s1_translator:av_readdata
	wire    [1:0] fft_in_0_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_0_s1_translator:av_address -> FFT_in_0:address
	wire   [31:0] fft_in_0_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_0:readdata -> FFT_in_0_s1_translator:av_readdata
	wire    [1:0] fft_in_1_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_1_s1_translator:av_address -> FFT_in_1:address
	wire   [31:0] fft_in_1_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_1:readdata -> FFT_in_1_s1_translator:av_readdata
	wire    [1:0] fft_in_2_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_2_s1_translator:av_address -> FFT_in_2:address
	wire   [31:0] fft_in_2_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_2:readdata -> FFT_in_2_s1_translator:av_readdata
	wire    [1:0] fft_in_3_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_3_s1_translator:av_address -> FFT_in_3:address
	wire   [31:0] fft_in_3_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_3:readdata -> FFT_in_3_s1_translator:av_readdata
	wire    [1:0] rotary_in_s1_translator_avalon_anti_slave_0_address;                                                                 // rotary_in_s1_translator:av_address -> rotary_in:address
	wire   [31:0] rotary_in_s1_translator_avalon_anti_slave_0_readdata;                                                                // rotary_in:readdata -> rotary_in_s1_translator:av_readdata
	wire    [1:0] fft_in_4_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_4_s1_translator:av_address -> FFT_in_4:address
	wire   [31:0] fft_in_4_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_4:readdata -> FFT_in_4_s1_translator:av_readdata
	wire    [1:0] fft_in_5_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_5_s1_translator:av_address -> FFT_in_5:address
	wire   [31:0] fft_in_5_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_5:readdata -> FFT_in_5_s1_translator:av_readdata
	wire    [1:0] fft_in_6_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_6_s1_translator:av_address -> FFT_in_6:address
	wire   [31:0] fft_in_6_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_6:readdata -> FFT_in_6_s1_translator:av_readdata
	wire    [1:0] fft_in_7_s1_translator_avalon_anti_slave_0_address;                                                                  // FFT_in_7_s1_translator:av_address -> FFT_in_7:address
	wire   [31:0] fft_in_7_s1_translator_avalon_anti_slave_0_readdata;                                                                 // FFT_in_7:readdata -> FFT_in_7_s1_translator:av_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                              // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                               // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                                 // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                                    // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                                   // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                                    // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                                // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                             // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                              // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                           // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest;                           // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_waitrequest
	wire    [1:0] vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount;                            // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_burstcount -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata;                             // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_writedata -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_address;                               // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_address -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock;                                  // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_lock -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_write;                                 // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_write -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_read;                                  // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_read -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata;                              // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_readdata
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess;                           // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_debugaccess -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable;                            // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_byteenable -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid;                         // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                                    // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                                     // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                                      // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                                        // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                                           // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                                          // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                                           // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                                       // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                                    // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                                     // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                                  // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // SRAM_avalon_sram_slave_translator:uav_waitrequest -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SRAM_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SRAM_avalon_sram_slave_translator:uav_writedata
	wire   [31:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                                         // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> SRAM_avalon_sram_slave_translator:uav_address
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                                           // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> SRAM_avalon_sram_slave_translator:uav_write
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                            // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SRAM_avalon_sram_slave_translator:uav_lock
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                                            // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> SRAM_avalon_sram_slave_translator:uav_read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // SRAM_avalon_sram_slave_translator:uav_readdata -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // SRAM_avalon_sram_slave_translator:uav_readdatavalid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SRAM_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SRAM_avalon_sram_slave_translator:uav_byteenable
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	wire    [3:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                      // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                             // red_led_pio_s1_translator:uav_waitrequest -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                              // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> red_led_pio_s1_translator:uav_burstcount
	wire   [31:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                               // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> red_led_pio_s1_translator:uav_writedata
	wire   [31:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                 // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> red_led_pio_s1_translator:uav_address
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                   // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> red_led_pio_s1_translator:uav_write
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                    // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> red_led_pio_s1_translator:uav_lock
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                    // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> red_led_pio_s1_translator:uav_read
	wire   [31:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                // red_led_pio_s1_translator:uav_readdata -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                           // red_led_pio_s1_translator:uav_readdatavalid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                             // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> red_led_pio_s1_translator:uav_debugaccess
	wire    [3:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                              // red_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> red_led_pio_s1_translator:uav_byteenable
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                      // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                            // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                    // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                             // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                            // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                   // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                         // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                 // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                          // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                         // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                       // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                        // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                       // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                       // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                        // red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                       // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // VGA_Character_buffer_avalon_char_control_slave_translator:uav_waitrequest -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_burstcount
	wire   [31:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_writedata
	wire   [31:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_address
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_write
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_lock
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_read
	wire   [31:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // VGA_Character_buffer_avalon_char_control_slave_translator:uav_readdata -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // VGA_Character_buffer_avalon_char_control_slave_translator:uav_readdatavalid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_debugaccess
	wire    [3:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Character_buffer_avalon_char_control_slave_translator:uav_byteenable
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_waitrequest -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_burstcount
	wire    [7:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_writedata
	wire   [31:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_address
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_write
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_lock
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_read
	wire    [7:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_readdata -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_readdatavalid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_debugaccess
	wire    [0:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Character_buffer_avalon_char_buffer_slave_translator:uav_byteenable
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire    [9:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;        // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;         // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;        // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // VGA_Pixel_Buffer_avalon_control_slave_translator:uav_waitrequest -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_burstcount
	wire   [31:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_writedata
	wire   [31:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_address
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_write
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_lock
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_read
	wire   [31:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // VGA_Pixel_Buffer_avalon_control_slave_translator:uav_readdata -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // VGA_Pixel_Buffer_avalon_control_slave_translator:uav_readdatavalid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_debugaccess
	wire    [3:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Pixel_Buffer_avalon_control_slave_translator:uav_byteenable
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // green_led_pio_s1_translator:uav_waitrequest -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> green_led_pio_s1_translator:uav_burstcount
	wire   [31:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> green_led_pio_s1_translator:uav_writedata
	wire   [31:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> green_led_pio_s1_translator:uav_address
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> green_led_pio_s1_translator:uav_write
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> green_led_pio_s1_translator:uav_lock
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> green_led_pio_s1_translator:uav_read
	wire   [31:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // green_led_pio_s1_translator:uav_readdata -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // green_led_pio_s1_translator:uav_readdatavalid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> green_led_pio_s1_translator:uav_debugaccess
	wire    [3:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // green_led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> green_led_pio_s1_translator:uav_byteenable
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                     // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                      // green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                     // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // control_in_s1_translator:uav_waitrequest -> control_in_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] control_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // control_in_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> control_in_s1_translator:uav_burstcount
	wire   [31:0] control_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // control_in_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> control_in_s1_translator:uav_writedata
	wire   [31:0] control_in_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                  // control_in_s1_translator_avalon_universal_slave_0_agent:m0_address -> control_in_s1_translator:uav_address
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                    // control_in_s1_translator_avalon_universal_slave_0_agent:m0_write -> control_in_s1_translator:uav_write
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // control_in_s1_translator_avalon_universal_slave_0_agent:m0_lock -> control_in_s1_translator:uav_lock
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                     // control_in_s1_translator_avalon_universal_slave_0_agent:m0_read -> control_in_s1_translator:uav_read
	wire   [31:0] control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // control_in_s1_translator:uav_readdata -> control_in_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // control_in_s1_translator:uav_readdatavalid -> control_in_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // control_in_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> control_in_s1_translator:uav_debugaccess
	wire    [3:0] control_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // control_in_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> control_in_s1_translator:uav_byteenable
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // control_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                        // control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                         // control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                        // control_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                             // control_out_s1_translator:uav_waitrequest -> control_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] control_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                              // control_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> control_out_s1_translator:uav_burstcount
	wire   [31:0] control_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                               // control_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> control_out_s1_translator:uav_writedata
	wire   [31:0] control_out_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                 // control_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> control_out_s1_translator:uav_address
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                   // control_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> control_out_s1_translator:uav_write
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                    // control_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> control_out_s1_translator:uav_lock
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                    // control_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> control_out_s1_translator:uav_read
	wire   [31:0] control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                // control_out_s1_translator:uav_readdata -> control_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                           // control_out_s1_translator:uav_readdatavalid -> control_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                             // control_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> control_out_s1_translator:uav_debugaccess
	wire    [3:0] control_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                              // control_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> control_out_s1_translator:uav_byteenable
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                      // control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                            // control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                    // control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                             // control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                            // control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                   // control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                         // control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                 // control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                          // control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                         // control_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                       // control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                        // control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                       // control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                       // control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                        // control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                       // control_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_0_s1_translator:uav_waitrequest -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_0_s1_translator:uav_burstcount
	wire   [31:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_0_s1_translator:uav_writedata
	wire   [31:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_0_s1_translator:uav_address
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_0_s1_translator:uav_write
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_0_s1_translator:uav_lock
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_0_s1_translator:uav_read
	wire   [31:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_0_s1_translator:uav_readdata -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_0_s1_translator:uav_readdatavalid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_0_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_0_s1_translator:uav_byteenable
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_1_s1_translator:uav_waitrequest -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_1_s1_translator:uav_burstcount
	wire   [31:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_1_s1_translator:uav_writedata
	wire   [31:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_1_s1_translator:uav_address
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_1_s1_translator:uav_write
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_1_s1_translator:uav_lock
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_1_s1_translator:uav_read
	wire   [31:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_1_s1_translator:uav_readdata -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_1_s1_translator:uav_readdatavalid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_1_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_1_s1_translator:uav_byteenable
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_2_s1_translator:uav_waitrequest -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_2_s1_translator:uav_burstcount
	wire   [31:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_2_s1_translator:uav_writedata
	wire   [31:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_2_s1_translator:uav_address
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_2_s1_translator:uav_write
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_2_s1_translator:uav_lock
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_2_s1_translator:uav_read
	wire   [31:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_2_s1_translator:uav_readdata -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_2_s1_translator:uav_readdatavalid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_2_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_2_s1_translator:uav_byteenable
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_3_s1_translator:uav_waitrequest -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_3_s1_translator:uav_burstcount
	wire   [31:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_3_s1_translator:uav_writedata
	wire   [31:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_3_s1_translator:uav_address
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_3_s1_translator:uav_write
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_3_s1_translator:uav_lock
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_3_s1_translator:uav_read
	wire   [31:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_3_s1_translator:uav_readdata -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_3_s1_translator:uav_readdatavalid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_3_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_3_s1_translator:uav_byteenable
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                               // rotary_in_s1_translator:uav_waitrequest -> rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> rotary_in_s1_translator:uav_burstcount
	wire   [31:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                 // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> rotary_in_s1_translator:uav_writedata
	wire   [31:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                   // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_address -> rotary_in_s1_translator:uav_address
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                     // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_write -> rotary_in_s1_translator:uav_write
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                      // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_lock -> rotary_in_s1_translator:uav_lock
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                      // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_read -> rotary_in_s1_translator:uav_read
	wire   [31:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                  // rotary_in_s1_translator:uav_readdata -> rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                             // rotary_in_s1_translator:uav_readdatavalid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                               // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rotary_in_s1_translator:uav_debugaccess
	wire    [3:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                // rotary_in_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> rotary_in_s1_translator:uav_byteenable
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                        // rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                              // rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                      // rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                               // rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                              // rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                     // rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                           // rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                   // rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                            // rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                           // rotary_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                         // rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                          // rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                         // rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                         // rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                          // rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                         // rotary_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_4_s1_translator:uav_waitrequest -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_4_s1_translator:uav_burstcount
	wire   [31:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_4_s1_translator:uav_writedata
	wire   [31:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_4_s1_translator:uav_address
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_4_s1_translator:uav_write
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_4_s1_translator:uav_lock
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_4_s1_translator:uav_read
	wire   [31:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_4_s1_translator:uav_readdata -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_4_s1_translator:uav_readdatavalid -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_4_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_4_s1_translator:uav_byteenable
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_5_s1_translator:uav_waitrequest -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_5_s1_translator:uav_burstcount
	wire   [31:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_5_s1_translator:uav_writedata
	wire   [31:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_5_s1_translator:uav_address
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_5_s1_translator:uav_write
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_5_s1_translator:uav_lock
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_5_s1_translator:uav_read
	wire   [31:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_5_s1_translator:uav_readdata -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_5_s1_translator:uav_readdatavalid -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_5_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_5_s1_translator:uav_byteenable
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_6_s1_translator:uav_waitrequest -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_6_s1_translator:uav_burstcount
	wire   [31:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_6_s1_translator:uav_writedata
	wire   [31:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_6_s1_translator:uav_address
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_6_s1_translator:uav_write
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_6_s1_translator:uav_lock
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_6_s1_translator:uav_read
	wire   [31:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_6_s1_translator:uav_readdata -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_6_s1_translator:uav_readdatavalid -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_6_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_6_s1_translator:uav_byteenable
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // FFT_in_7_s1_translator:uav_waitrequest -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FFT_in_7_s1_translator:uav_burstcount
	wire   [31:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FFT_in_7_s1_translator:uav_writedata
	wire   [31:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_address -> FFT_in_7_s1_translator:uav_address
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_write -> FFT_in_7_s1_translator:uav_write
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FFT_in_7_s1_translator:uav_lock
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_read -> FFT_in_7_s1_translator:uav_read
	wire   [31:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // FFT_in_7_s1_translator:uav_readdata -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // FFT_in_7_s1_translator:uav_readdatavalid -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FFT_in_7_s1_translator:uav_debugaccess
	wire    [3:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FFT_in_7_s1_translator:uav_byteenable
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                    // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                          // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                  // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [108:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                           // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                          // addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                        // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire   [90:0] vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data;                         // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                           // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                                 // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                         // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [108:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                                  // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                                 // addr_router_002:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [108:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                           // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [90:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                                            // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_001:sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [108:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [108:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_003:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [108:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_004:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                             // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                   // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                           // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [108:0] red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                    // red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                   // id_router_005:sink_ready -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [108:0] vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [81:0] vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_007:sink_ready -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [108:0] vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_008:sink_ready -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [108:0] green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_009:sink_ready -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // control_in_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // control_in_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // control_in_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [108:0] control_in_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                     // control_in_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          control_in_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_010:sink_ready -> control_in_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                             // control_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                   // control_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                           // control_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [108:0] control_out_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                    // control_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          control_out_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                   // id_router_011:sink_ready -> control_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [108:0] fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_012:sink_ready -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [108:0] fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_013:sink_ready -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [108:0] fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_014:sink_ready -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [108:0] fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_015:sink_ready -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                               // rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                     // rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                             // rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [108:0] rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                      // rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                     // id_router_016:sink_ready -> rotary_in_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [108:0] fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_017:sink_ready -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [108:0] fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_018:sink_ready -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [108:0] fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_019:sink_ready -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [108:0] fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_020:sink_ready -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                                   // burst_adapter:source0_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                         // burst_adapter:source0_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                                 // burst_adapter:source0_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] burst_adapter_source0_data;                                                                                          // burst_adapter:source0_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                         // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [20:0] burst_adapter_source0_channel;                                                                                       // burst_adapter:source0_channel -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                               // burst_adapter_001:source0_endofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                                     // burst_adapter_001:source0_valid -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                             // burst_adapter_001:source0_startofpacket -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] burst_adapter_001_source0_data;                                                                                      // burst_adapter_001:source0_data -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                                     // VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [20:0] burst_adapter_001_source0_channel;                                                                                   // burst_adapter_001:source0_channel -> VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                      // rst_controller:reset_out -> [addr_router:reset, addr_router_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:in_reset, crosser_007:out_reset, crosser_008:out_reset, crosser_009:out_reset, id_router:reset, id_router_002:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_002:reset, rsp_xbar_mux:reset, rsp_xbar_mux_002:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset]
	wire          external_clocks_sys_clk_reset_reset;                                                                                 // external_clocks:sys_reset_n -> rst_controller:reset_in1
	wire          rst_controller_001_reset_out_reset;                                                                                  // rst_controller_001:reset_out -> [FFT_in_0:reset_n, FFT_in_0_s1_translator:reset, FFT_in_0_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_1:reset_n, FFT_in_1_s1_translator:reset, FFT_in_1_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_2:reset_n, FFT_in_2_s1_translator:reset, FFT_in_2_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_3:reset_n, FFT_in_3_s1_translator:reset, FFT_in_3_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_4:reset_n, FFT_in_4_s1_translator:reset, FFT_in_4_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_5:reset_n, FFT_in_5_s1_translator:reset, FFT_in_5_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_6:reset_n, FFT_in_6_s1_translator:reset, FFT_in_6_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FFT_in_7:reset_n, FFT_in_7_s1_translator:reset, FFT_in_7_s1_translator_avalon_universal_slave_0_agent:reset, FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FFT_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, control_in:reset_n, control_in_s1_translator:reset, control_in_s1_translator_avalon_universal_slave_0_agent:reset, control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, control_out:reset_n, control_out_s1_translator:reset, control_out_s1_translator_avalon_universal_slave_0_agent:reset, control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, external_clocks:reset, green_led_pio:reset_n, green_led_pio_s1_translator:reset, green_led_pio_s1_translator_avalon_universal_slave_0_agent:reset, green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, red_led_pio:reset_n, red_led_pio_s1_translator:reset, red_led_pio_s1_translator_avalon_universal_slave_0_agent:reset, red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rotary_in:reset_n, rotary_in_s1_translator:reset, rotary_in_s1_translator_avalon_universal_slave_0_agent:reset, rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, sys_clk_timer:reset_n, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_002_reset_out_reset;                                                                                  // rst_controller_002:reset_out -> [Alpha_Blending:reset, SRAM:reset, SRAM_avalon_sram_slave_translator:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Character_buffer:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, VGA_Character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Character_buffer_avalon_char_control_slave_translator:reset, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Dual_Clock_FIFO:reset_stream_in, VGA_Pixel_Buffer:reset, VGA_Pixel_Buffer_avalon_control_slave_translator:reset, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator:reset, VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, VGA_Scaler:reset, VGA_pixel_RGB_Resampler:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux_001:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:in_reset, crosser_008:in_reset, crosser_009:in_reset, id_router_001:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset]
	wire          cpu_jtag_debug_module_reset_reset;                                                                                   // cpu:jtag_debug_module_resetrequest -> [rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire          rst_controller_003_reset_out_reset;                                                                                  // rst_controller_003:reset_out -> [VGA_Controller:reset, VGA_Dual_Clock_FIFO:reset_stream_out]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src0_data;                                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [20:0] cmd_xbar_demux_src0_channel;                                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [90:0] cmd_xbar_demux_001_src0_data;                                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_001:sink1_data
	wire   [20:0] cmd_xbar_demux_001_src0_channel;                                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                                 // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                       // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                               // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src0_data;                                                                                        // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux:sink1_data
	wire   [20:0] cmd_xbar_demux_002_src0_channel;                                                                                     // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                                                 // cmd_xbar_demux_002:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                                       // cmd_xbar_demux_002:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                                               // cmd_xbar_demux_002:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src2_data;                                                                                        // cmd_xbar_demux_002:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src2_channel;                                                                                     // cmd_xbar_demux_002:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src3_endofpacket;                                                                                 // cmd_xbar_demux_002:src3_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src3_valid;                                                                                       // cmd_xbar_demux_002:src3_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src3_startofpacket;                                                                               // cmd_xbar_demux_002:src3_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src3_data;                                                                                        // cmd_xbar_demux_002:src3_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src3_channel;                                                                                     // cmd_xbar_demux_002:src3_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src4_endofpacket;                                                                                 // cmd_xbar_demux_002:src4_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src4_valid;                                                                                       // cmd_xbar_demux_002:src4_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src4_startofpacket;                                                                               // cmd_xbar_demux_002:src4_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src4_data;                                                                                        // cmd_xbar_demux_002:src4_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src4_channel;                                                                                     // cmd_xbar_demux_002:src4_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src5_endofpacket;                                                                                 // cmd_xbar_demux_002:src5_endofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src5_valid;                                                                                       // cmd_xbar_demux_002:src5_valid -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src5_startofpacket;                                                                               // cmd_xbar_demux_002:src5_startofpacket -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src5_data;                                                                                        // cmd_xbar_demux_002:src5_data -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src5_channel;                                                                                     // cmd_xbar_demux_002:src5_channel -> red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src9_endofpacket;                                                                                 // cmd_xbar_demux_002:src9_endofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src9_valid;                                                                                       // cmd_xbar_demux_002:src9_valid -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src9_startofpacket;                                                                               // cmd_xbar_demux_002:src9_startofpacket -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src9_data;                                                                                        // cmd_xbar_demux_002:src9_data -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src9_channel;                                                                                     // cmd_xbar_demux_002:src9_channel -> green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src10_endofpacket;                                                                                // cmd_xbar_demux_002:src10_endofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src10_valid;                                                                                      // cmd_xbar_demux_002:src10_valid -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src10_startofpacket;                                                                              // cmd_xbar_demux_002:src10_startofpacket -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src10_data;                                                                                       // cmd_xbar_demux_002:src10_data -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src10_channel;                                                                                    // cmd_xbar_demux_002:src10_channel -> control_in_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src11_endofpacket;                                                                                // cmd_xbar_demux_002:src11_endofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src11_valid;                                                                                      // cmd_xbar_demux_002:src11_valid -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src11_startofpacket;                                                                              // cmd_xbar_demux_002:src11_startofpacket -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src11_data;                                                                                       // cmd_xbar_demux_002:src11_data -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src11_channel;                                                                                    // cmd_xbar_demux_002:src11_channel -> control_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src12_endofpacket;                                                                                // cmd_xbar_demux_002:src12_endofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src12_valid;                                                                                      // cmd_xbar_demux_002:src12_valid -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src12_startofpacket;                                                                              // cmd_xbar_demux_002:src12_startofpacket -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src12_data;                                                                                       // cmd_xbar_demux_002:src12_data -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src12_channel;                                                                                    // cmd_xbar_demux_002:src12_channel -> FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src13_endofpacket;                                                                                // cmd_xbar_demux_002:src13_endofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src13_valid;                                                                                      // cmd_xbar_demux_002:src13_valid -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src13_startofpacket;                                                                              // cmd_xbar_demux_002:src13_startofpacket -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src13_data;                                                                                       // cmd_xbar_demux_002:src13_data -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src13_channel;                                                                                    // cmd_xbar_demux_002:src13_channel -> FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src14_endofpacket;                                                                                // cmd_xbar_demux_002:src14_endofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src14_valid;                                                                                      // cmd_xbar_demux_002:src14_valid -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src14_startofpacket;                                                                              // cmd_xbar_demux_002:src14_startofpacket -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src14_data;                                                                                       // cmd_xbar_demux_002:src14_data -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src14_channel;                                                                                    // cmd_xbar_demux_002:src14_channel -> FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src15_endofpacket;                                                                                // cmd_xbar_demux_002:src15_endofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src15_valid;                                                                                      // cmd_xbar_demux_002:src15_valid -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src15_startofpacket;                                                                              // cmd_xbar_demux_002:src15_startofpacket -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src15_data;                                                                                       // cmd_xbar_demux_002:src15_data -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src15_channel;                                                                                    // cmd_xbar_demux_002:src15_channel -> FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src16_endofpacket;                                                                                // cmd_xbar_demux_002:src16_endofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src16_valid;                                                                                      // cmd_xbar_demux_002:src16_valid -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src16_startofpacket;                                                                              // cmd_xbar_demux_002:src16_startofpacket -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src16_data;                                                                                       // cmd_xbar_demux_002:src16_data -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src16_channel;                                                                                    // cmd_xbar_demux_002:src16_channel -> rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src17_endofpacket;                                                                                // cmd_xbar_demux_002:src17_endofpacket -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src17_valid;                                                                                      // cmd_xbar_demux_002:src17_valid -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src17_startofpacket;                                                                              // cmd_xbar_demux_002:src17_startofpacket -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src17_data;                                                                                       // cmd_xbar_demux_002:src17_data -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src17_channel;                                                                                    // cmd_xbar_demux_002:src17_channel -> FFT_in_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src18_endofpacket;                                                                                // cmd_xbar_demux_002:src18_endofpacket -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src18_valid;                                                                                      // cmd_xbar_demux_002:src18_valid -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src18_startofpacket;                                                                              // cmd_xbar_demux_002:src18_startofpacket -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src18_data;                                                                                       // cmd_xbar_demux_002:src18_data -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src18_channel;                                                                                    // cmd_xbar_demux_002:src18_channel -> FFT_in_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src19_endofpacket;                                                                                // cmd_xbar_demux_002:src19_endofpacket -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src19_valid;                                                                                      // cmd_xbar_demux_002:src19_valid -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src19_startofpacket;                                                                              // cmd_xbar_demux_002:src19_startofpacket -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src19_data;                                                                                       // cmd_xbar_demux_002:src19_data -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src19_channel;                                                                                    // cmd_xbar_demux_002:src19_channel -> FFT_in_6_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src20_endofpacket;                                                                                // cmd_xbar_demux_002:src20_endofpacket -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src20_valid;                                                                                      // cmd_xbar_demux_002:src20_valid -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src20_startofpacket;                                                                              // cmd_xbar_demux_002:src20_startofpacket -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src20_data;                                                                                       // cmd_xbar_demux_002:src20_data -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_demux_002_src20_channel;                                                                                    // cmd_xbar_demux_002:src20_channel -> FFT_in_7_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [108:0] rsp_xbar_demux_src0_data;                                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [20:0] rsp_xbar_demux_src0_channel;                                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [108:0] rsp_xbar_demux_src1_data;                                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_002:sink0_data
	wire   [20:0] rsp_xbar_demux_src1_channel;                                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                           // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                                 // rsp_xbar_demux_001:src1_endofpacket -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                       // rsp_xbar_demux_001:src1_valid -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                               // rsp_xbar_demux_001:src1_startofpacket -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [90:0] rsp_xbar_demux_001_src1_data;                                                                                        // rsp_xbar_demux_001:src1_data -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [20:0] rsp_xbar_demux_001_src1_channel;                                                                                     // rsp_xbar_demux_001:src1_channel -> VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [108:0] rsp_xbar_demux_002_src0_data;                                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_002:sink2_data
	wire   [20:0] rsp_xbar_demux_002_src0_channel;                                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                       // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_002:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [108:0] rsp_xbar_demux_003_src0_data;                                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_002:sink3_data
	wire   [20:0] rsp_xbar_demux_003_src0_channel;                                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_002:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                       // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                                 // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                       // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_002:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                               // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [108:0] rsp_xbar_demux_004_src0_data;                                                                                        // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_002:sink4_data
	wire   [20:0] rsp_xbar_demux_004_src0_channel;                                                                                     // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_002:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                       // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_002:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	wire  [108:0] rsp_xbar_demux_005_src0_data;                                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_002:sink5_data
	wire   [20:0] rsp_xbar_demux_005_src0_channel;                                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_002:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                       // rsp_xbar_mux_002:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                                 // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_002:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                       // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_002:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                               // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_002:sink9_startofpacket
	wire  [108:0] rsp_xbar_demux_009_src0_data;                                                                                        // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_002:sink9_data
	wire   [20:0] rsp_xbar_demux_009_src0_channel;                                                                                     // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_002:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                       // rsp_xbar_mux_002:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                                 // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_002:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                       // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_002:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                               // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_002:sink10_startofpacket
	wire  [108:0] rsp_xbar_demux_010_src0_data;                                                                                        // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_002:sink10_data
	wire   [20:0] rsp_xbar_demux_010_src0_channel;                                                                                     // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_002:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                       // rsp_xbar_mux_002:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                                 // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_002:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                       // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_002:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                               // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_002:sink11_startofpacket
	wire  [108:0] rsp_xbar_demux_011_src0_data;                                                                                        // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_002:sink11_data
	wire   [20:0] rsp_xbar_demux_011_src0_channel;                                                                                     // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_002:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                       // rsp_xbar_mux_002:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                                 // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_002:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                       // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_002:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                               // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_002:sink12_startofpacket
	wire  [108:0] rsp_xbar_demux_012_src0_data;                                                                                        // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_002:sink12_data
	wire   [20:0] rsp_xbar_demux_012_src0_channel;                                                                                     // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_002:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                       // rsp_xbar_mux_002:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                                 // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_002:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                       // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_002:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                               // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_002:sink13_startofpacket
	wire  [108:0] rsp_xbar_demux_013_src0_data;                                                                                        // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_002:sink13_data
	wire   [20:0] rsp_xbar_demux_013_src0_channel;                                                                                     // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_002:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                       // rsp_xbar_mux_002:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                                 // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_002:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                       // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_002:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                               // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_002:sink14_startofpacket
	wire  [108:0] rsp_xbar_demux_014_src0_data;                                                                                        // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_002:sink14_data
	wire   [20:0] rsp_xbar_demux_014_src0_channel;                                                                                     // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_002:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                       // rsp_xbar_mux_002:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                                 // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_002:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                       // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_002:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                               // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_002:sink15_startofpacket
	wire  [108:0] rsp_xbar_demux_015_src0_data;                                                                                        // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_002:sink15_data
	wire   [20:0] rsp_xbar_demux_015_src0_channel;                                                                                     // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_002:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                       // rsp_xbar_mux_002:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                                 // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_002:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                       // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_002:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                               // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_002:sink16_startofpacket
	wire  [108:0] rsp_xbar_demux_016_src0_data;                                                                                        // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_002:sink16_data
	wire   [20:0] rsp_xbar_demux_016_src0_channel;                                                                                     // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_002:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                       // rsp_xbar_mux_002:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                                 // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_002:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                       // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_002:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                               // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_002:sink17_startofpacket
	wire  [108:0] rsp_xbar_demux_017_src0_data;                                                                                        // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_002:sink17_data
	wire   [20:0] rsp_xbar_demux_017_src0_channel;                                                                                     // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_002:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                       // rsp_xbar_mux_002:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                                 // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_002:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                       // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_002:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                               // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_002:sink18_startofpacket
	wire  [108:0] rsp_xbar_demux_018_src0_data;                                                                                        // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_002:sink18_data
	wire   [20:0] rsp_xbar_demux_018_src0_channel;                                                                                     // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_002:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                       // rsp_xbar_mux_002:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                                 // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_002:sink19_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                                       // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_002:sink19_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                               // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_002:sink19_startofpacket
	wire  [108:0] rsp_xbar_demux_019_src0_data;                                                                                        // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_002:sink19_data
	wire   [20:0] rsp_xbar_demux_019_src0_channel;                                                                                     // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_002:sink19_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                                       // rsp_xbar_mux_002:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                                 // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_002:sink20_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                                       // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_002:sink20_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                                               // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_002:sink20_startofpacket
	wire  [108:0] rsp_xbar_demux_020_src0_data;                                                                                        // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_002:sink20_data
	wire   [20:0] rsp_xbar_demux_020_src0_channel;                                                                                     // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_002:sink20_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                                       // rsp_xbar_mux_002:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire          addr_router_src_endofpacket;                                                                                         // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                               // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                                       // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [108:0] addr_router_src_data;                                                                                                // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [20:0] addr_router_src_channel;                                                                                             // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                               // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                        // rsp_xbar_mux:src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                              // rsp_xbar_mux:src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                      // rsp_xbar_mux:src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] rsp_xbar_mux_src_data;                                                                                               // rsp_xbar_mux:src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [20:0] rsp_xbar_mux_src_channel;                                                                                            // rsp_xbar_mux:src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                                     // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                           // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                                   // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire   [90:0] addr_router_001_src_data;                                                                                            // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [20:0] addr_router_001_src_channel;                                                                                         // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                           // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_demux_001_src1_ready;                                                                                       // VGA_Pixel_Buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src1_ready
	wire          addr_router_002_src_endofpacket;                                                                                     // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                           // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                                   // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [108:0] addr_router_002_src_data;                                                                                            // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [20:0] addr_router_002_src_channel;                                                                                         // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                           // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                                    // rsp_xbar_mux_002:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                                          // rsp_xbar_mux_002:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                                  // rsp_xbar_mux_002:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] rsp_xbar_mux_002_src_data;                                                                                           // rsp_xbar_mux_002:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [20:0] rsp_xbar_mux_002_src_channel;                                                                                        // rsp_xbar_mux_002:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                                          // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                        // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                              // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                      // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_src_data;                                                                                               // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] cmd_xbar_mux_src_channel;                                                                                            // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [108:0] id_router_src_data;                                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [20:0] id_router_src_channel;                                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                                    // cmd_xbar_mux_001:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                          // cmd_xbar_mux_001:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                                  // cmd_xbar_mux_001:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [90:0] cmd_xbar_mux_001_src_data;                                                                                           // cmd_xbar_mux_001:src_data -> burst_adapter:sink0_data
	wire   [20:0] cmd_xbar_mux_001_src_channel;                                                                                        // cmd_xbar_mux_001:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                          // burst_adapter:sink0_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                       // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                             // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                     // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [90:0] id_router_001_src_data;                                                                                              // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [20:0] id_router_001_src_channel;                                                                                           // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                             // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_002_src2_ready;                                                                                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src2_ready
	wire          id_router_002_src_endofpacket;                                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [108:0] id_router_002_src_data;                                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [20:0] id_router_002_src_channel;                                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_002_src3_ready;                                                                                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src3_ready
	wire          id_router_003_src_endofpacket;                                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [108:0] id_router_003_src_data;                                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [20:0] id_router_003_src_channel;                                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_002_src4_ready;                                                                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [108:0] id_router_004_src_data;                                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [20:0] id_router_004_src_channel;                                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_002_src5_ready;                                                                                       // red_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src5_ready
	wire          id_router_005_src_endofpacket;                                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [108:0] id_router_005_src_data;                                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [20:0] id_router_005_src_channel;                                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          crosser_out_ready;                                                                                                   // VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_006_src_endofpacket;                                                                                       // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                             // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                     // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [108:0] id_router_006_src_data;                                                                                              // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [20:0] id_router_006_src_channel;                                                                                           // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                             // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          crosser_006_out_ready;                                                                                               // burst_adapter_001:sink0_ready -> crosser_006:out_ready
	wire          id_router_007_src_endofpacket;                                                                                       // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                             // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                     // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [81:0] id_router_007_src_data;                                                                                              // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [20:0] id_router_007_src_channel;                                                                                           // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                             // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          crosser_001_out_ready;                                                                                               // VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire          id_router_008_src_endofpacket;                                                                                       // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                             // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                     // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [108:0] id_router_008_src_data;                                                                                              // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [20:0] id_router_008_src_channel;                                                                                           // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                             // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_002_src9_ready;                                                                                       // green_led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src9_ready
	wire          id_router_009_src_endofpacket;                                                                                       // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                             // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                     // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [108:0] id_router_009_src_data;                                                                                              // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [20:0] id_router_009_src_channel;                                                                                           // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                             // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_002_src10_ready;                                                                                      // control_in_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src10_ready
	wire          id_router_010_src_endofpacket;                                                                                       // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                             // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                     // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [108:0] id_router_010_src_data;                                                                                              // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [20:0] id_router_010_src_channel;                                                                                           // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                             // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_002_src11_ready;                                                                                      // control_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src11_ready
	wire          id_router_011_src_endofpacket;                                                                                       // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                             // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                     // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [108:0] id_router_011_src_data;                                                                                              // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [20:0] id_router_011_src_channel;                                                                                           // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                             // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_002_src12_ready;                                                                                      // FFT_in_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src12_ready
	wire          id_router_012_src_endofpacket;                                                                                       // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                             // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                     // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [108:0] id_router_012_src_data;                                                                                              // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [20:0] id_router_012_src_channel;                                                                                           // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                             // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_002_src13_ready;                                                                                      // FFT_in_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src13_ready
	wire          id_router_013_src_endofpacket;                                                                                       // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                             // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                     // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [108:0] id_router_013_src_data;                                                                                              // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [20:0] id_router_013_src_channel;                                                                                           // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                             // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_002_src14_ready;                                                                                      // FFT_in_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src14_ready
	wire          id_router_014_src_endofpacket;                                                                                       // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                             // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                     // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [108:0] id_router_014_src_data;                                                                                              // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [20:0] id_router_014_src_channel;                                                                                           // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                             // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_002_src15_ready;                                                                                      // FFT_in_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src15_ready
	wire          id_router_015_src_endofpacket;                                                                                       // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                             // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                     // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [108:0] id_router_015_src_data;                                                                                              // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [20:0] id_router_015_src_channel;                                                                                           // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                             // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_002_src16_ready;                                                                                      // rotary_in_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src16_ready
	wire          id_router_016_src_endofpacket;                                                                                       // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                             // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                     // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [108:0] id_router_016_src_data;                                                                                              // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [20:0] id_router_016_src_channel;                                                                                           // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                             // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_002_src17_ready;                                                                                      // FFT_in_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src17_ready
	wire          id_router_017_src_endofpacket;                                                                                       // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                             // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                     // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [108:0] id_router_017_src_data;                                                                                              // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [20:0] id_router_017_src_channel;                                                                                           // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                             // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_002_src18_ready;                                                                                      // FFT_in_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src18_ready
	wire          id_router_018_src_endofpacket;                                                                                       // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                             // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                     // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [108:0] id_router_018_src_data;                                                                                              // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [20:0] id_router_018_src_channel;                                                                                           // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                             // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_002_src19_ready;                                                                                      // FFT_in_6_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src19_ready
	wire          id_router_019_src_endofpacket;                                                                                       // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                                             // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                                     // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [108:0] id_router_019_src_data;                                                                                              // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [20:0] id_router_019_src_channel;                                                                                           // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                                             // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_002_src20_ready;                                                                                      // FFT_in_7_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src20_ready
	wire          id_router_020_src_endofpacket;                                                                                       // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                                             // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                                     // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [108:0] id_router_020_src_data;                                                                                              // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [20:0] id_router_020_src_channel;                                                                                           // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                                             // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                     // cmd_xbar_demux:src1_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                           // cmd_xbar_demux:src1_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                                   // cmd_xbar_demux:src1_startofpacket -> width_adapter:in_startofpacket
	wire  [108:0] cmd_xbar_demux_src1_data;                                                                                            // cmd_xbar_demux:src1_data -> width_adapter:in_data
	wire   [20:0] cmd_xbar_demux_src1_channel;                                                                                         // cmd_xbar_demux:src1_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                           // width_adapter:in_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                                 // cmd_xbar_demux_002:src1_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                                       // cmd_xbar_demux_002:src1_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                                               // cmd_xbar_demux_002:src1_startofpacket -> width_adapter_001:in_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src1_data;                                                                                        // cmd_xbar_demux_002:src1_data -> width_adapter_001:in_data
	wire   [20:0] cmd_xbar_demux_002_src1_channel;                                                                                     // cmd_xbar_demux_002:src1_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                                       // width_adapter_001:in_ready -> cmd_xbar_demux_002:src1_ready
	wire          cmd_xbar_demux_002_src7_endofpacket;                                                                                 // cmd_xbar_demux_002:src7_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_002_src7_valid;                                                                                       // cmd_xbar_demux_002:src7_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_002_src7_startofpacket;                                                                               // cmd_xbar_demux_002:src7_startofpacket -> width_adapter_002:in_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src7_data;                                                                                        // cmd_xbar_demux_002:src7_data -> width_adapter_002:in_data
	wire   [20:0] cmd_xbar_demux_002_src7_channel;                                                                                     // cmd_xbar_demux_002:src7_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_002_src7_ready;                                                                                       // width_adapter_002:in_ready -> cmd_xbar_demux_002:src7_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                                 // rsp_xbar_demux_001:src0_endofpacket -> width_adapter_003:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                       // rsp_xbar_demux_001:src0_valid -> width_adapter_003:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                               // rsp_xbar_demux_001:src0_startofpacket -> width_adapter_003:in_startofpacket
	wire   [90:0] rsp_xbar_demux_001_src0_data;                                                                                        // rsp_xbar_demux_001:src0_data -> width_adapter_003:in_data
	wire   [20:0] rsp_xbar_demux_001_src0_channel;                                                                                     // rsp_xbar_demux_001:src0_channel -> width_adapter_003:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                       // width_adapter_003:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                                                 // rsp_xbar_demux_001:src2_endofpacket -> width_adapter_004:in_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                                       // rsp_xbar_demux_001:src2_valid -> width_adapter_004:in_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                                               // rsp_xbar_demux_001:src2_startofpacket -> width_adapter_004:in_startofpacket
	wire   [90:0] rsp_xbar_demux_001_src2_data;                                                                                        // rsp_xbar_demux_001:src2_data -> width_adapter_004:in_data
	wire   [20:0] rsp_xbar_demux_001_src2_channel;                                                                                     // rsp_xbar_demux_001:src2_channel -> width_adapter_004:in_channel
	wire          rsp_xbar_demux_001_src2_ready;                                                                                       // width_adapter_004:in_ready -> rsp_xbar_demux_001:src2_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                                 // rsp_xbar_demux_007:src0_endofpacket -> width_adapter_005:in_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                       // rsp_xbar_demux_007:src0_valid -> width_adapter_005:in_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                               // rsp_xbar_demux_007:src0_startofpacket -> width_adapter_005:in_startofpacket
	wire   [81:0] rsp_xbar_demux_007_src0_data;                                                                                        // rsp_xbar_demux_007:src0_data -> width_adapter_005:in_data
	wire   [20:0] rsp_xbar_demux_007_src0_channel;                                                                                     // rsp_xbar_demux_007:src0_channel -> width_adapter_005:in_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                       // width_adapter_005:in_ready -> rsp_xbar_demux_007:src0_ready
	wire          crosser_out_endofpacket;                                                                                             // crosser:out_endofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                                   // crosser:out_valid -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                                           // crosser:out_startofpacket -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] crosser_out_data;                                                                                                    // crosser:out_data -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] crosser_out_channel;                                                                                                 // crosser:out_channel -> VGA_Character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src6_endofpacket;                                                                                 // cmd_xbar_demux_002:src6_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_002_src6_valid;                                                                                       // cmd_xbar_demux_002:src6_valid -> crosser:in_valid
	wire          cmd_xbar_demux_002_src6_startofpacket;                                                                               // cmd_xbar_demux_002:src6_startofpacket -> crosser:in_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src6_data;                                                                                        // cmd_xbar_demux_002:src6_data -> crosser:in_data
	wire   [20:0] cmd_xbar_demux_002_src6_channel;                                                                                     // cmd_xbar_demux_002:src6_channel -> crosser:in_channel
	wire          cmd_xbar_demux_002_src6_ready;                                                                                       // crosser:in_ready -> cmd_xbar_demux_002:src6_ready
	wire          crosser_001_out_endofpacket;                                                                                         // crosser_001:out_endofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_001_out_valid;                                                                                               // crosser_001:out_valid -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_001_out_startofpacket;                                                                                       // crosser_001:out_startofpacket -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] crosser_001_out_data;                                                                                                // crosser_001:out_data -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [20:0] crosser_001_out_channel;                                                                                             // crosser_001:out_channel -> VGA_Pixel_Buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src8_endofpacket;                                                                                 // cmd_xbar_demux_002:src8_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_002_src8_valid;                                                                                       // cmd_xbar_demux_002:src8_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_002_src8_startofpacket;                                                                               // cmd_xbar_demux_002:src8_startofpacket -> crosser_001:in_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src8_data;                                                                                        // cmd_xbar_demux_002:src8_data -> crosser_001:in_data
	wire   [20:0] cmd_xbar_demux_002_src8_channel;                                                                                     // cmd_xbar_demux_002:src8_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_002_src8_ready;                                                                                       // crosser_001:in_ready -> cmd_xbar_demux_002:src8_ready
	wire          crosser_002_out_endofpacket;                                                                                         // crosser_002:out_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	wire          crosser_002_out_valid;                                                                                               // crosser_002:out_valid -> rsp_xbar_mux_002:sink6_valid
	wire          crosser_002_out_startofpacket;                                                                                       // crosser_002:out_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	wire  [108:0] crosser_002_out_data;                                                                                                // crosser_002:out_data -> rsp_xbar_mux_002:sink6_data
	wire   [20:0] crosser_002_out_channel;                                                                                             // crosser_002:out_channel -> rsp_xbar_mux_002:sink6_channel
	wire          crosser_002_out_ready;                                                                                               // rsp_xbar_mux_002:sink6_ready -> crosser_002:out_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                                 // rsp_xbar_demux_006:src0_endofpacket -> crosser_002:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                       // rsp_xbar_demux_006:src0_valid -> crosser_002:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                               // rsp_xbar_demux_006:src0_startofpacket -> crosser_002:in_startofpacket
	wire  [108:0] rsp_xbar_demux_006_src0_data;                                                                                        // rsp_xbar_demux_006:src0_data -> crosser_002:in_data
	wire   [20:0] rsp_xbar_demux_006_src0_channel;                                                                                     // rsp_xbar_demux_006:src0_channel -> crosser_002:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                       // crosser_002:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          crosser_003_out_endofpacket;                                                                                         // crosser_003:out_endofpacket -> rsp_xbar_mux_002:sink8_endofpacket
	wire          crosser_003_out_valid;                                                                                               // crosser_003:out_valid -> rsp_xbar_mux_002:sink8_valid
	wire          crosser_003_out_startofpacket;                                                                                       // crosser_003:out_startofpacket -> rsp_xbar_mux_002:sink8_startofpacket
	wire  [108:0] crosser_003_out_data;                                                                                                // crosser_003:out_data -> rsp_xbar_mux_002:sink8_data
	wire   [20:0] crosser_003_out_channel;                                                                                             // crosser_003:out_channel -> rsp_xbar_mux_002:sink8_channel
	wire          crosser_003_out_ready;                                                                                               // rsp_xbar_mux_002:sink8_ready -> crosser_003:out_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                                 // rsp_xbar_demux_008:src0_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                       // rsp_xbar_demux_008:src0_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                               // rsp_xbar_demux_008:src0_startofpacket -> crosser_003:in_startofpacket
	wire  [108:0] rsp_xbar_demux_008_src0_data;                                                                                        // rsp_xbar_demux_008:src0_data -> crosser_003:in_data
	wire   [20:0] rsp_xbar_demux_008_src0_channel;                                                                                     // rsp_xbar_demux_008:src0_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                       // crosser_003:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          crosser_004_out_endofpacket;                                                                                         // crosser_004:out_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          crosser_004_out_valid;                                                                                               // crosser_004:out_valid -> cmd_xbar_mux_001:sink0_valid
	wire          crosser_004_out_startofpacket;                                                                                       // crosser_004:out_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [90:0] crosser_004_out_data;                                                                                                // crosser_004:out_data -> cmd_xbar_mux_001:sink0_data
	wire   [20:0] crosser_004_out_channel;                                                                                             // crosser_004:out_channel -> cmd_xbar_mux_001:sink0_channel
	wire          crosser_004_out_ready;                                                                                               // cmd_xbar_mux_001:sink0_ready -> crosser_004:out_ready
	wire          width_adapter_src_endofpacket;                                                                                       // width_adapter:out_endofpacket -> crosser_004:in_endofpacket
	wire          width_adapter_src_valid;                                                                                             // width_adapter:out_valid -> crosser_004:in_valid
	wire          width_adapter_src_startofpacket;                                                                                     // width_adapter:out_startofpacket -> crosser_004:in_startofpacket
	wire   [90:0] width_adapter_src_data;                                                                                              // width_adapter:out_data -> crosser_004:in_data
	wire          width_adapter_src_ready;                                                                                             // crosser_004:in_ready -> width_adapter:out_ready
	wire   [20:0] width_adapter_src_channel;                                                                                           // width_adapter:out_channel -> crosser_004:in_channel
	wire          crosser_005_out_endofpacket;                                                                                         // crosser_005:out_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          crosser_005_out_valid;                                                                                               // crosser_005:out_valid -> cmd_xbar_mux_001:sink2_valid
	wire          crosser_005_out_startofpacket;                                                                                       // crosser_005:out_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire   [90:0] crosser_005_out_data;                                                                                                // crosser_005:out_data -> cmd_xbar_mux_001:sink2_data
	wire   [20:0] crosser_005_out_channel;                                                                                             // crosser_005:out_channel -> cmd_xbar_mux_001:sink2_channel
	wire          crosser_005_out_ready;                                                                                               // cmd_xbar_mux_001:sink2_ready -> crosser_005:out_ready
	wire          width_adapter_001_src_endofpacket;                                                                                   // width_adapter_001:out_endofpacket -> crosser_005:in_endofpacket
	wire          width_adapter_001_src_valid;                                                                                         // width_adapter_001:out_valid -> crosser_005:in_valid
	wire          width_adapter_001_src_startofpacket;                                                                                 // width_adapter_001:out_startofpacket -> crosser_005:in_startofpacket
	wire   [90:0] width_adapter_001_src_data;                                                                                          // width_adapter_001:out_data -> crosser_005:in_data
	wire          width_adapter_001_src_ready;                                                                                         // crosser_005:in_ready -> width_adapter_001:out_ready
	wire   [20:0] width_adapter_001_src_channel;                                                                                       // width_adapter_001:out_channel -> crosser_005:in_channel
	wire          crosser_006_out_endofpacket;                                                                                         // crosser_006:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          crosser_006_out_valid;                                                                                               // crosser_006:out_valid -> burst_adapter_001:sink0_valid
	wire          crosser_006_out_startofpacket;                                                                                       // crosser_006:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [81:0] crosser_006_out_data;                                                                                                // crosser_006:out_data -> burst_adapter_001:sink0_data
	wire   [20:0] crosser_006_out_channel;                                                                                             // crosser_006:out_channel -> burst_adapter_001:sink0_channel
	wire          width_adapter_002_src_endofpacket;                                                                                   // width_adapter_002:out_endofpacket -> crosser_006:in_endofpacket
	wire          width_adapter_002_src_valid;                                                                                         // width_adapter_002:out_valid -> crosser_006:in_valid
	wire          width_adapter_002_src_startofpacket;                                                                                 // width_adapter_002:out_startofpacket -> crosser_006:in_startofpacket
	wire   [81:0] width_adapter_002_src_data;                                                                                          // width_adapter_002:out_data -> crosser_006:in_data
	wire          width_adapter_002_src_ready;                                                                                         // crosser_006:in_ready -> width_adapter_002:out_ready
	wire   [20:0] width_adapter_002_src_channel;                                                                                       // width_adapter_002:out_channel -> crosser_006:in_channel
	wire          crosser_007_out_endofpacket;                                                                                         // crosser_007:out_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          crosser_007_out_valid;                                                                                               // crosser_007:out_valid -> rsp_xbar_mux:sink1_valid
	wire          crosser_007_out_startofpacket;                                                                                       // crosser_007:out_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [108:0] crosser_007_out_data;                                                                                                // crosser_007:out_data -> rsp_xbar_mux:sink1_data
	wire   [20:0] crosser_007_out_channel;                                                                                             // crosser_007:out_channel -> rsp_xbar_mux:sink1_channel
	wire          crosser_007_out_ready;                                                                                               // rsp_xbar_mux:sink1_ready -> crosser_007:out_ready
	wire          width_adapter_003_src_endofpacket;                                                                                   // width_adapter_003:out_endofpacket -> crosser_007:in_endofpacket
	wire          width_adapter_003_src_valid;                                                                                         // width_adapter_003:out_valid -> crosser_007:in_valid
	wire          width_adapter_003_src_startofpacket;                                                                                 // width_adapter_003:out_startofpacket -> crosser_007:in_startofpacket
	wire  [108:0] width_adapter_003_src_data;                                                                                          // width_adapter_003:out_data -> crosser_007:in_data
	wire          width_adapter_003_src_ready;                                                                                         // crosser_007:in_ready -> width_adapter_003:out_ready
	wire   [20:0] width_adapter_003_src_channel;                                                                                       // width_adapter_003:out_channel -> crosser_007:in_channel
	wire          crosser_008_out_endofpacket;                                                                                         // crosser_008:out_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          crosser_008_out_valid;                                                                                               // crosser_008:out_valid -> rsp_xbar_mux_002:sink1_valid
	wire          crosser_008_out_startofpacket;                                                                                       // crosser_008:out_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [108:0] crosser_008_out_data;                                                                                                // crosser_008:out_data -> rsp_xbar_mux_002:sink1_data
	wire   [20:0] crosser_008_out_channel;                                                                                             // crosser_008:out_channel -> rsp_xbar_mux_002:sink1_channel
	wire          crosser_008_out_ready;                                                                                               // rsp_xbar_mux_002:sink1_ready -> crosser_008:out_ready
	wire          width_adapter_004_src_endofpacket;                                                                                   // width_adapter_004:out_endofpacket -> crosser_008:in_endofpacket
	wire          width_adapter_004_src_valid;                                                                                         // width_adapter_004:out_valid -> crosser_008:in_valid
	wire          width_adapter_004_src_startofpacket;                                                                                 // width_adapter_004:out_startofpacket -> crosser_008:in_startofpacket
	wire  [108:0] width_adapter_004_src_data;                                                                                          // width_adapter_004:out_data -> crosser_008:in_data
	wire          width_adapter_004_src_ready;                                                                                         // crosser_008:in_ready -> width_adapter_004:out_ready
	wire   [20:0] width_adapter_004_src_channel;                                                                                       // width_adapter_004:out_channel -> crosser_008:in_channel
	wire          crosser_009_out_endofpacket;                                                                                         // crosser_009:out_endofpacket -> rsp_xbar_mux_002:sink7_endofpacket
	wire          crosser_009_out_valid;                                                                                               // crosser_009:out_valid -> rsp_xbar_mux_002:sink7_valid
	wire          crosser_009_out_startofpacket;                                                                                       // crosser_009:out_startofpacket -> rsp_xbar_mux_002:sink7_startofpacket
	wire  [108:0] crosser_009_out_data;                                                                                                // crosser_009:out_data -> rsp_xbar_mux_002:sink7_data
	wire   [20:0] crosser_009_out_channel;                                                                                             // crosser_009:out_channel -> rsp_xbar_mux_002:sink7_channel
	wire          crosser_009_out_ready;                                                                                               // rsp_xbar_mux_002:sink7_ready -> crosser_009:out_ready
	wire          width_adapter_005_src_endofpacket;                                                                                   // width_adapter_005:out_endofpacket -> crosser_009:in_endofpacket
	wire          width_adapter_005_src_valid;                                                                                         // width_adapter_005:out_valid -> crosser_009:in_valid
	wire          width_adapter_005_src_startofpacket;                                                                                 // width_adapter_005:out_startofpacket -> crosser_009:in_startofpacket
	wire  [108:0] width_adapter_005_src_data;                                                                                          // width_adapter_005:out_data -> crosser_009:in_data
	wire          width_adapter_005_src_ready;                                                                                         // crosser_009:in_ready -> width_adapter_005:out_ready
	wire   [20:0] width_adapter_005_src_channel;                                                                                       // width_adapter_005:out_channel -> crosser_009:in_channel
	wire          irq_mapper_receiver0_irq;                                                                                            // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                            // sys_clk_timer:irq -> irq_mapper:receiver1_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                                       // irq_mapper:sender_irq -> cpu:d_irq

	nios2VGA_cpu cpu (
		.clk                                   (clk_clk),                                                          //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                  // custom_instruction_master.readra
	);

	nios2VGA_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	nios2VGA_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                                    //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        // reset.reset_n
		.address    (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_clk_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                                    //   irq.irq
	);

	nios2VGA_sysid sysid (
		.clock    (clk_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	nios2VGA_red_led_pio red_led_pio (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (red_led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~red_led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (red_led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (red_led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (red_led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (red_led_pio_external_connection_export)                    // external_connection.export
	);

	nios2VGA_external_clocks external_clocks (
		.CLOCK_50    (clk_clk),                             //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset),  // clk_in_primary_reset.reset
		.sys_clk     (external_clocks_sys_clk_clk),         //              sys_clk.clk
		.sys_reset_n (external_clocks_sys_clk_reset_reset), //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clock_clk),                     //            sdram_clk.clk
		.VGA_CLK     (vga_clock_out_clk_clk)                //              vga_clk.clk
	);

	nios2VGA_VGA_Dual_Clock_FIFO vga_dual_clock_fifo (
		.clk_stream_in            (external_clocks_sys_clk_clk),                               //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_002_reset_out_reset),                        //   clock_stream_in_reset.reset
		.clk_stream_out           (vga_clock_out_clk_clk),                                     //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_003_reset_out_reset),                        //  clock_stream_out_reset.reset
		.stream_in_ready          (alpha_blending_avalon_blended_source_ready),                //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (alpha_blending_avalon_blended_source_startofpacket),        //                        .startofpacket
		.stream_in_endofpacket    (alpha_blending_avalon_blended_source_endofpacket),          //                        .endofpacket
		.stream_in_valid          (alpha_blending_avalon_blended_source_valid),                //                        .valid
		.stream_in_data           (alpha_blending_avalon_blended_source_data),                 //                        .data
		.stream_out_ready         (vga_dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (vga_dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (vga_dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	nios2VGA_Alpha_Blending alpha_blending (
		.clk                      (external_clocks_sys_clk_clk),                           //            clock_reset.clk
		.reset                    (rst_controller_002_reset_out_reset),                    //      clock_reset_reset.reset
		.foreground_data          (vga_character_buffer_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (vga_character_buffer_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (vga_character_buffer_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (vga_character_buffer_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (vga_character_buffer_avalon_char_source_ready),         //                       .ready
		.background_data          (vga_scaler_avalon_scaler_source_data),                  // avalon_background_sink.data
		.background_startofpacket (vga_scaler_avalon_scaler_source_startofpacket),         //                       .startofpacket
		.background_endofpacket   (vga_scaler_avalon_scaler_source_endofpacket),           //                       .endofpacket
		.background_valid         (vga_scaler_avalon_scaler_source_valid),                 //                       .valid
		.background_ready         (vga_scaler_avalon_scaler_source_ready),                 //                       .ready
		.output_ready             (alpha_blending_avalon_blended_source_ready),            //  avalon_blended_source.ready
		.output_data              (alpha_blending_avalon_blended_source_data),             //                       .data
		.output_startofpacket     (alpha_blending_avalon_blended_source_startofpacket),    //                       .startofpacket
		.output_endofpacket       (alpha_blending_avalon_blended_source_endofpacket),      //                       .endofpacket
		.output_valid             (alpha_blending_avalon_blended_source_valid)             //                       .valid
	);

	nios2VGA_VGA_Controller vga_controller (
		.clk           (vga_clock_out_clk_clk),                                     //        clock_reset.clk
		.reset         (rst_controller_003_reset_out_reset),                        //  clock_reset_reset.reset
		.data          (vga_dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (vga_dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (vga_dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_external_CLK),                               // external_interface.export
		.VGA_HS        (vga_controller_external_HS),                                //                   .export
		.VGA_VS        (vga_controller_external_VS),                                //                   .export
		.VGA_BLANK     (vga_controller_external_BLANK),                             //                   .export
		.VGA_SYNC      (vga_controller_external_SYNC),                              //                   .export
		.VGA_R         (vga_controller_external_R),                                 //                   .export
		.VGA_G         (vga_controller_external_G),                                 //                   .export
		.VGA_B         (vga_controller_external_B)                                  //                   .export
	);

	nios2VGA_VGA_Character_buffer vga_character_buffer (
		.clk                  (external_clocks_sys_clk_clk),                                                              //               clock_reset.clk
		.reset                (rst_controller_002_reset_out_reset),                                                       //         clock_reset_reset.reset
		.ctrl_address         (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable), //                          .byteenable
		.ctrl_chipselect      (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect), //                          .chipselect
		.ctrl_read            (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),       //                          .read
		.ctrl_write           (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),      //                          .write
		.ctrl_writedata       (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),  //                          .writedata
		.ctrl_readdata        (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),   //                          .readdata
		.buf_byteenable       (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),  //                          .chipselect
		.buf_read             (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),        //                          .read
		.buf_write            (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),       //                          .write
		.buf_writedata        (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.buf_readdata         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.buf_waitrequest      (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.buf_address          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),     //                          .address
		.stream_ready         (vga_character_buffer_avalon_char_source_ready),                                            //        avalon_char_source.ready
		.stream_startofpacket (vga_character_buffer_avalon_char_source_startofpacket),                                    //                          .startofpacket
		.stream_endofpacket   (vga_character_buffer_avalon_char_source_endofpacket),                                      //                          .endofpacket
		.stream_valid         (vga_character_buffer_avalon_char_source_valid),                                            //                          .valid
		.stream_data          (vga_character_buffer_avalon_char_source_data)                                              //                          .data
	);

	nios2VGA_VGA_Scaler vga_scaler (
		.clk                      (external_clocks_sys_clk_clk),                             //          clock_reset.clk
		.reset                    (rst_controller_002_reset_out_reset),                      //    clock_reset_reset.reset
		.stream_in_startofpacket  (vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (vga_pixel_rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (vga_pixel_rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (vga_pixel_rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (vga_scaler_avalon_scaler_source_ready),                   // avalon_scaler_source.ready
		.stream_out_startofpacket (vga_scaler_avalon_scaler_source_startofpacket),           //                     .startofpacket
		.stream_out_endofpacket   (vga_scaler_avalon_scaler_source_endofpacket),             //                     .endofpacket
		.stream_out_valid         (vga_scaler_avalon_scaler_source_valid),                   //                     .valid
		.stream_out_data          (vga_scaler_avalon_scaler_source_data)                     //                     .data
	);

	nios2VGA_VGA_pixel_RGB_Resampler vga_pixel_rgb_resampler (
		.clk                      (external_clocks_sys_clk_clk),                             //       clock_reset.clk
		.reset                    (rst_controller_002_reset_out_reset),                      // clock_reset_reset.reset
		.stream_in_startofpacket  (vga_pixel_buffer_avalon_pixel_source_startofpacket),      //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (vga_pixel_buffer_avalon_pixel_source_endofpacket),        //                  .endofpacket
		.stream_in_valid          (vga_pixel_buffer_avalon_pixel_source_valid),              //                  .valid
		.stream_in_ready          (vga_pixel_buffer_avalon_pixel_source_ready),              //                  .ready
		.stream_in_data           (vga_pixel_buffer_avalon_pixel_source_data),               //                  .data
		.stream_out_ready         (vga_pixel_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (vga_pixel_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (vga_pixel_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	nios2VGA_VGA_Pixel_Buffer vga_pixel_buffer (
		.clk                  (external_clocks_sys_clk_clk),                                                     //             clock_reset.clk
		.reset                (rst_controller_002_reset_out_reset),                                              //       clock_reset_reset.reset
		.master_readdatavalid (vga_pixel_buffer_avalon_pixel_dma_master_readdatavalid),                          // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (vga_pixel_buffer_avalon_pixel_dma_master_waitrequest),                            //                        .waitrequest
		.master_address       (vga_pixel_buffer_avalon_pixel_dma_master_address),                                //                        .address
		.master_arbiterlock   (vga_pixel_buffer_avalon_pixel_dma_master_lock),                                   //                        .lock
		.master_read          (vga_pixel_buffer_avalon_pixel_dma_master_read),                                   //                        .read
		.master_readdata      (vga_pixel_buffer_avalon_pixel_dma_master_readdata),                               //                        .readdata
		.slave_address        (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_address),    //    avalon_control_slave.address
		.slave_byteenable     (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_byteenable), //                        .byteenable
		.slave_read           (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_read),       //                        .read
		.slave_write          (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_write),      //                        .write
		.slave_writedata      (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_writedata),  //                        .writedata
		.slave_readdata       (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_readdata),   //                        .readdata
		.stream_ready         (vga_pixel_buffer_avalon_pixel_source_ready),                                      //     avalon_pixel_source.ready
		.stream_startofpacket (vga_pixel_buffer_avalon_pixel_source_startofpacket),                              //                        .startofpacket
		.stream_endofpacket   (vga_pixel_buffer_avalon_pixel_source_endofpacket),                                //                        .endofpacket
		.stream_valid         (vga_pixel_buffer_avalon_pixel_source_valid),                                      //                        .valid
		.stream_data          (vga_pixel_buffer_avalon_pixel_source_data)                                        //                        .data
	);

	nios2VGA_SRAM sram (
		.clk           (external_clocks_sys_clk_clk),                                         //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),                                  //  clock_reset_reset.reset
		.SRAM_DQ       (sram_external_interface_DQ),                                          // external_interface.export
		.SRAM_ADDR     (sram_external_interface_ADDR),                                        //                   .export
		.SRAM_LB_N     (sram_external_interface_LB_N),                                        //                   .export
		.SRAM_UB_N     (sram_external_interface_UB_N),                                        //                   .export
		.SRAM_CE_N     (sram_external_interface_CE_N),                                        //                   .export
		.SRAM_OE_N     (sram_external_interface_OE_N),                                        //                   .export
		.SRAM_WE_N     (sram_external_interface_WE_N),                                        //                   .export
		.address       (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	nios2VGA_green_led_pio green_led_pio (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (green_led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~green_led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (green_led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (green_led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (green_led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (green_led_pio_external_connection_export)                    // external_connection.export
	);

	nios2VGA_control_in control_in (
		.clk      (clk_clk),                                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address  (control_in_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (control_in_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (nios_cntrl_in_export)                                   // external_connection.export
	);

	nios2VGA_control_out control_out (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (control_out_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~control_out_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (control_out_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (control_out_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (control_out_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (nios_cntrl_out_export)                                     // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_0 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_0_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_0_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_0_export)                                      // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_1 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_1_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_1_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_1_export)                                      // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_2 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_2_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_2_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_2_export)                                      // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_3 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_3_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_3_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_3_export)                                      // external_connection.export
	);

	nios2VGA_control_in rotary_in (
		.clk      (clk_clk),                                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address  (rotary_in_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (rotary_in_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (rotary_in_export)                                      // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_4 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_4_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_4_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_4_export)                                      // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_5 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_5_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_5_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_5_export)                                      // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_6 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_6_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_6_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_6_export)                                      // external_connection.export
	);

	nios2VGA_FFT_in_0 fft_in_7 (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (fft_in_7_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (fft_in_7_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (fft_in_7_export)                                      // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                      (clk_clk),                                                                   //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_byteenable            (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                          //               (terminated)
		.av_write                 (1'b0),                                                                      //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) vga_pixel_buffer_avalon_pixel_dma_master_translator (
		.clk                      (external_clocks_sys_clk_clk),                                                                 //                       clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                          //                     reset.reset
		.uav_address              (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (vga_pixel_buffer_avalon_pixel_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (vga_pixel_buffer_avalon_pixel_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (vga_pixel_buffer_avalon_pixel_dma_master_read),                                               //                          .read
		.av_readdata              (vga_pixel_buffer_avalon_pixel_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (vga_pixel_buffer_avalon_pixel_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock                  (vga_pixel_buffer_avalon_pixel_dma_master_lock),                                               //                          .lock
		.av_burstcount            (1'b1),                                                                                        //               (terminated)
		.av_byteenable            (2'b11),                                                                                       //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                                        //               (terminated)
		.av_write                 (1'b0),                                                                                        //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                                        //               (terminated)
		.uav_clken                (),                                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                                       //               (terminated)
		.av_response              (),                                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_data_master_translator (
		.clk                      (clk_clk),                                                            //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address              (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_data_master_read),                                               //                          .read
		.av_readdata              (cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_data_master_write),                                              //                          .write
		.av_writedata             (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_readdatavalid         (),                                                                   //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_avalon_sram_slave_translator (
		.clk                      (external_clocks_sys_clk_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                //                    reset.reset
		.uav_address              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_chipselect            (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_clk_timer_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sys_clk_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) red_led_pio_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (red_led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (red_led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (red_led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (red_led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (red_led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) vga_character_buffer_avalon_char_control_slave_translator (
		.clk                      (external_clocks_sys_clk_clk),                                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                                        //                    reset.reset
		.uav_address              (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (vga_character_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                                          //              (terminated)
		.av_lock                  (),                                                                                                          //              (terminated)
		.av_clken                 (),                                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                                          //              (terminated)
		.uav_response             (),                                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) vga_character_buffer_avalon_char_buffer_slave_translator (
		.clk                      (external_clocks_sys_clk_clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                                       //                    reset.reset
		.uav_address              (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                                         //              (terminated)
		.av_lock                  (),                                                                                                         //              (terminated)
		.av_clken                 (),                                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                                         //              (terminated)
		.uav_response             (),                                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) vga_pixel_buffer_avalon_control_slave_translator (
		.clk                      (external_clocks_sys_clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                               //                    reset.reset
		.uav_address              (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (vga_pixel_buffer_avalon_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                                 //              (terminated)
		.av_lock                  (),                                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                                 //              (terminated)
		.av_clken                 (),                                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                                 //              (terminated)
		.uav_response             (),                                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) green_led_pio_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (green_led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (green_led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (green_led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (green_led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (green_led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) control_in_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (control_in_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (control_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (control_in_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (control_in_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (control_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (control_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (control_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (control_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (control_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (control_in_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (control_in_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                         //              (terminated)
		.av_read                  (),                                                                         //              (terminated)
		.av_writedata             (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_chipselect            (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) control_out_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (control_out_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (control_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (control_out_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (control_out_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (control_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (control_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (control_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (control_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (control_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (control_out_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (control_out_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (control_out_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (control_out_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (control_out_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_0_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_1_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_2_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_3_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rotary_in_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (rotary_in_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (rotary_in_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_writedata             (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_chipselect            (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_4_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_5_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_6_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_6_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_6_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fft_in_7_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fft_in_7_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (fft_in_7_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (21),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                            //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                             //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                              //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                           //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                       //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                             //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (81),
		.PKT_THREAD_ID_L           (81),
		.PKT_CACHE_H               (88),
		.PKT_CACHE_L               (85),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (21),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (external_clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                   // clk_reset.reset
		.av_address              (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_001_src1_valid),                                                                        //        rp.valid
		.rp_data                 (rsp_xbar_demux_001_src1_data),                                                                         //          .data
		.rp_channel              (rsp_xbar_demux_001_src1_channel),                                                                      //          .channel
		.rp_startofpacket        (rsp_xbar_demux_001_src1_startofpacket),                                                                //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_001_src1_endofpacket),                                                                  //          .endofpacket
		.rp_ready                (rsp_xbar_demux_001_src1_ready),                                                                        //          .ready
		.av_response             (),                                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (21),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                     //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address              (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_002_src_valid),                                                  //        rp.valid
		.rp_data                 (rsp_xbar_mux_002_src_data),                                                   //          .data
		.rp_channel              (rsp_xbar_mux_002_src_channel),                                                //          .channel
		.rp_startofpacket        (rsp_xbar_mux_002_src_startofpacket),                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_002_src_endofpacket),                                            //          .endofpacket
		.rp_ready                (rsp_xbar_mux_002_src_ready),                                                  //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_startofpacket  (1'b0),                                                                                 // (terminated)
		.in_endofpacket    (1'b0),                                                                                 // (terminated)
		.out_startofpacket (),                                                                                     // (terminated)
		.out_endofpacket   (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (external_clocks_sys_clk_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                 //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                 //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                  //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                           //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                               //                .channel
		.rf_sink_ready           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src2_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src2_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_002_src2_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src2_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src2_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src2_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src3_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src3_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_002_src3_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src3_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src3_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src3_channel),                                                       //                .channel
		.rf_sink_ready           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src4_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src4_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_002_src4_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src4_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src4_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src4_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_startofpacket  (1'b0),                                                                               // (terminated)
		.in_endofpacket    (1'b0),                                                                               // (terminated)
		.out_startofpacket (),                                                                                   // (terminated)
		.out_endofpacket   (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) red_led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (red_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src5_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src5_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_002_src5_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src5_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src5_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src5_channel),                                                     //                .channel
		.rf_sink_ready           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                          // (terminated)
		.out_startofpacket (),                                                                              // (terminated)
		.out_endofpacket   (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (external_clocks_sys_clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                                  //       clk_reset.reset
		.m0_address              (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                                                   //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                                                   //                .valid
		.cp_data                 (crosser_out_data),                                                                                                    //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                                                           //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                                             //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                                                 //                .channel
		.rf_sink_ready           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                                  // clk_reset.reset
		.in_data           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                // (terminated)
		.almost_full_data  (),                                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                                // (terminated)
		.out_empty         (),                                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                                // (terminated)
		.out_error         (),                                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                                // (terminated)
		.out_channel       ()                                                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                          // (terminated)
		.almost_full_data  (),                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                                                          // (terminated)
		.out_startofpacket (),                                                                                                              // (terminated)
		.out_endofpacket   (),                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                          // (terminated)
		.out_empty         (),                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                          // (terminated)
		.out_error         (),                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                          // (terminated)
		.out_channel       ()                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (66),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (67),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (external_clocks_sys_clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                                 //       clk_reset.reset
		.m0_address              (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                                    //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                                    //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                                     //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                                              //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                                  //                .channel
		.rf_sink_ready           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                                 // clk_reset.reset
		.in_data           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                               // (terminated)
		.almost_full_data  (),                                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                                               // (terminated)
		.out_empty         (),                                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                                               // (terminated)
		.out_error         (),                                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                                               // (terminated)
		.out_channel       ()                                                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (10),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                           // clk_reset.reset
		.in_data           (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                                         // (terminated)
		.csr_readdata      (),                                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                         // (terminated)
		.almost_full_data  (),                                                                                                             // (terminated)
		.almost_empty_data (),                                                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                                                         // (terminated)
		.out_startofpacket (),                                                                                                             // (terminated)
		.out_endofpacket   (),                                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                                         // (terminated)
		.out_empty         (),                                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                                         // (terminated)
		.out_error         (),                                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                                         // (terminated)
		.out_channel       ()                                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (external_clocks_sys_clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                                                      //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                                                      //                .valid
		.cp_data                 (crosser_001_out_data),                                                                                       //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                                              //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                                                //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                                                    //                .channel
		.rf_sink_ready           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (external_clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                                 // (terminated)
		.csr_readdata      (),                                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                 // (terminated)
		.almost_full_data  (),                                                                                                     // (terminated)
		.almost_empty_data (),                                                                                                     // (terminated)
		.in_startofpacket  (1'b0),                                                                                                 // (terminated)
		.in_endofpacket    (1'b0),                                                                                                 // (terminated)
		.out_startofpacket (),                                                                                                     // (terminated)
		.out_endofpacket   (),                                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                                 // (terminated)
		.out_empty         (),                                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                                 // (terminated)
		.out_error         (),                                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                                 // (terminated)
		.out_channel       ()                                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) green_led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (green_led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src9_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src9_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_002_src9_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src9_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src9_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src9_channel),                                                       //                .channel
		.rf_sink_ready           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) control_in_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (control_in_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (control_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (control_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (control_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (control_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (control_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (control_in_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (control_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (control_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (control_in_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (control_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (control_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (control_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (control_in_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (control_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src10_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src10_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_002_src10_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src10_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src10_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src10_channel),                                                   //                .channel
		.rf_sink_ready           (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (control_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (control_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (control_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) control_out_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (control_out_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (control_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (control_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (control_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (control_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (control_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (control_out_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (control_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (control_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (control_out_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (control_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (control_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (control_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (control_out_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (control_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src11_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src11_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_002_src11_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src11_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src11_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src11_channel),                                                    //                .channel
		.rf_sink_ready           (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (control_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (control_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (control_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                          // (terminated)
		.out_startofpacket (),                                                                              // (terminated)
		.out_endofpacket   (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src12_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src12_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src12_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src12_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src12_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src12_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src13_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src13_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src13_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src13_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src13_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src13_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src14_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src14_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src14_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src14_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src14_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src14_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src15_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src15_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src15_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src15_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src15_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src15_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rotary_in_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rotary_in_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src16_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src16_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_002_src16_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src16_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src16_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src16_channel),                                                  //                .channel
		.rf_sink_ready           (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rotary_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rotary_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src17_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src17_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src17_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src17_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src17_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src17_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src18_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src18_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src18_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src18_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src18_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src18_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_6_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_6_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src19_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src19_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src19_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src19_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src19_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src19_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (21),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fft_in_7_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fft_in_7_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src20_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src20_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_002_src20_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src20_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src20_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src20_channel),                                                 //                .channel
		.rf_sink_ready           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	nios2VGA_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios2VGA_addr_router_001 addr_router_001 (
		.sink_ready         (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_pixel_buffer_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (external_clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                                       //          .endofpacket
	);

	nios2VGA_addr_router_002 addr_router_002 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                   //          .valid
		.src_data           (addr_router_002_src_data),                                                    //          .data
		.src_channel        (addr_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                              //          .endofpacket
	);

	nios2VGA_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios2VGA_id_router_001 id_router_001 (
		.sink_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (external_clocks_sys_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                           //       src.ready
		.src_valid          (id_router_001_src_valid),                                                           //          .valid
		.src_data           (id_router_001_src_data),                                                            //          .data
		.src_channel        (id_router_001_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                      //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_002 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                //          .valid
		.src_data           (id_router_002_src_data),                                                                 //          .data
		.src_channel        (id_router_002_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_003 (
		.sink_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                     //       src.ready
		.src_valid          (id_router_003_src_valid),                                                     //          .valid
		.src_data           (id_router_003_src_data),                                                      //          .data
		.src_channel        (id_router_003_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_004 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                        //       src.ready
		.src_valid          (id_router_004_src_valid),                                                        //          .valid
		.src_data           (id_router_004_src_data),                                                         //          .data
		.src_channel        (id_router_004_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                   //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_005 (
		.sink_ready         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (red_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                   //       src.ready
		.src_valid          (id_router_005_src_valid),                                                   //          .valid
		.src_data           (id_router_005_src_data),                                                    //          .data
		.src_channel        (id_router_005_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                              //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_006 (
		.sink_ready         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_character_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (external_clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                                        // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                                   //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                                   //          .valid
		.src_data           (id_router_006_src_data),                                                                                    //          .data
		.src_channel        (id_router_006_src_channel),                                                                                 //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                           //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                              //          .endofpacket
	);

	nios2VGA_id_router_007 id_router_007 (
		.sink_ready         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_character_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (external_clocks_sys_clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                                  //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                                  //          .valid
		.src_data           (id_router_007_src_data),                                                                                   //          .data
		.src_channel        (id_router_007_src_channel),                                                                                //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                                          //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                                             //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_008 (
		.sink_ready         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_pixel_buffer_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (external_clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                          //          .valid
		.src_data           (id_router_008_src_data),                                                                           //          .data
		.src_channel        (id_router_008_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                     //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_009 (
		.sink_ready         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (green_led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                     //       src.ready
		.src_valid          (id_router_009_src_valid),                                                     //          .valid
		.src_data           (id_router_009_src_data),                                                      //          .data
		.src_channel        (id_router_009_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_010 (
		.sink_ready         (control_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (control_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (control_in_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (control_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (control_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                  //       src.ready
		.src_valid          (id_router_010_src_valid),                                                  //          .valid
		.src_data           (id_router_010_src_data),                                                   //          .data
		.src_channel        (id_router_010_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                             //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_011 (
		.sink_ready         (control_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (control_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (control_out_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (control_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (control_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                   //       src.ready
		.src_valid          (id_router_011_src_valid),                                                   //          .valid
		.src_data           (id_router_011_src_data),                                                    //          .data
		.src_channel        (id_router_011_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                              //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_012 (
		.sink_ready         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                //       src.ready
		.src_valid          (id_router_012_src_valid),                                                //          .valid
		.src_data           (id_router_012_src_data),                                                 //          .data
		.src_channel        (id_router_012_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_013 (
		.sink_ready         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                //       src.ready
		.src_valid          (id_router_013_src_valid),                                                //          .valid
		.src_data           (id_router_013_src_data),                                                 //          .data
		.src_channel        (id_router_013_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_014 (
		.sink_ready         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                //       src.ready
		.src_valid          (id_router_014_src_valid),                                                //          .valid
		.src_data           (id_router_014_src_data),                                                 //          .data
		.src_channel        (id_router_014_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_015 (
		.sink_ready         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                //       src.ready
		.src_valid          (id_router_015_src_valid),                                                //          .valid
		.src_data           (id_router_015_src_data),                                                 //          .data
		.src_channel        (id_router_015_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_016 (
		.sink_ready         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rotary_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                 //       src.ready
		.src_valid          (id_router_016_src_valid),                                                 //          .valid
		.src_data           (id_router_016_src_data),                                                  //          .data
		.src_channel        (id_router_016_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                            //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_017 (
		.sink_ready         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                //       src.ready
		.src_valid          (id_router_017_src_valid),                                                //          .valid
		.src_data           (id_router_017_src_data),                                                 //          .data
		.src_channel        (id_router_017_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_018 (
		.sink_ready         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                //       src.ready
		.src_valid          (id_router_018_src_valid),                                                //          .valid
		.src_data           (id_router_018_src_data),                                                 //          .data
		.src_channel        (id_router_018_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_019 (
		.sink_ready         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                //       src.ready
		.src_valid          (id_router_019_src_valid),                                                //          .valid
		.src_data           (id_router_019_src_data),                                                 //          .data
		.src_channel        (id_router_019_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                           //          .endofpacket
	);

	nios2VGA_id_router_002 id_router_020 (
		.sink_ready         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fft_in_7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                //       src.ready
		.src_valid          (id_router_020_src_valid),                                                //          .valid
		.src_data           (id_router_020_src_data),                                                 //          .data
		.src_channel        (id_router_020_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                           //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (21),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (external_clocks_sys_clk_clk),         //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_001_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_001_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_001_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_001_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_001_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_001_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (21),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (external_clocks_sys_clk_clk),             //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (crosser_006_out_valid),                   //     sink0.valid
		.sink0_data            (crosser_006_out_data),                    //          .data
		.sink0_channel         (crosser_006_out_channel),                 //          .channel
		.sink0_startofpacket   (crosser_006_out_startofpacket),           //          .startofpacket
		.sink0_endofpacket     (crosser_006_out_endofpacket),             //          .endofpacket
		.sink0_ready           (crosser_006_out_ready),                   //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                       // reset_in0.reset
		.reset_in1  (~external_clocks_sys_clk_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                              //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req  (),                                     // (terminated)
		.reset_in2  (1'b0),                                 // (terminated)
		.reset_in3  (1'b0),                                 // (terminated)
		.reset_in4  (1'b0),                                 // (terminated)
		.reset_in5  (1'b0),                                 // (terminated)
		.reset_in6  (1'b0),                                 // (terminated)
		.reset_in7  (1'b0),                                 // (terminated)
		.reset_in8  (1'b0),                                 // (terminated)
		.reset_in9  (1'b0),                                 // (terminated)
		.reset_in10 (1'b0),                                 // (terminated)
		.reset_in11 (1'b0),                                 // (terminated)
		.reset_in12 (1'b0),                                 // (terminated)
		.reset_in13 (1'b0),                                 // (terminated)
		.reset_in14 (1'b0),                                 // (terminated)
		.reset_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (external_clocks_sys_clk_clk),        //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (vga_clock_out_clk_clk),              //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios2VGA_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios2VGA_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (external_clocks_sys_clk_clk),           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_002_src_ready),              //      sink.ready
		.sink_channel        (addr_router_002_src_channel),            //          .channel
		.sink_data           (addr_router_002_src_data),               //          .data
		.sink_startofpacket  (addr_router_002_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_002_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_002_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_002_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_002_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_002_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_002_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_002_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_002_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_002_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_002_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_002_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_002_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_002_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_002_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_002_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_002_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_002_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_002_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_002_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_002_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_002_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_002_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_002_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_002_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_002_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_002_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_002_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_002_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_002_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_002_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_002_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_002_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_002_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_002_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_002_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_002_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_002_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_002_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_002_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_002_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_002_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_002_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_002_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_002_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_002_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_002_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_002_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_002_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_002_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_002_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_002_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_002_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_002_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_002_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_002_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_002_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_002_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_002_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_002_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_002_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_002_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_002_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_002_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_002_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_002_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_002_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_002_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_002_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_002_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_002_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_002_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_002_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_002_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_002_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_002_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_002_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_002_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_002_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_002_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_002_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_002_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_002_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_002_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_002_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_002_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_002_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_002_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_002_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_002_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_002_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_002_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_002_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_002_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_002_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_002_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_002_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_002_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_002_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_002_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_002_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_002_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_002_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_002_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_002_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_002_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_002_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_002_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_002_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_002_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_002_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_002_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_002_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_002_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_002_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_002_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_002_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_002_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_002_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_002_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_002_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_002_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_002_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_002_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_002_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_002_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_002_src20_endofpacket)    //          .endofpacket
	);

	nios2VGA_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (external_clocks_sys_clk_clk),           //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (crosser_004_out_ready),                 //     sink0.ready
		.sink0_valid         (crosser_004_out_valid),                 //          .valid
		.sink0_channel       (crosser_004_out_channel),               //          .channel
		.sink0_data          (crosser_004_out_data),                  //          .data
		.sink0_startofpacket (crosser_004_out_startofpacket),         //          .startofpacket
		.sink0_endofpacket   (crosser_004_out_endofpacket),           //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (crosser_005_out_ready),                 //     sink2.ready
		.sink2_valid         (crosser_005_out_valid),                 //          .valid
		.sink2_channel       (crosser_005_out_channel),               //          .channel
		.sink2_data          (crosser_005_out_data),                  //          .data
		.sink2_startofpacket (crosser_005_out_startofpacket),         //          .startofpacket
		.sink2_endofpacket   (crosser_005_out_endofpacket)            //          .endofpacket
	);

	nios2VGA_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (external_clocks_sys_clk_clk),           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (external_clocks_sys_clk_clk),           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_007 rsp_xbar_demux_007 (
		.clk                (external_clocks_sys_clk_clk),           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (external_clocks_sys_clk_clk),           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_018 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_demux_002 rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	nios2VGA_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                           //       clk.clk
		.reset               (rst_controller_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_007_out_ready),             //     sink1.ready
		.sink1_valid         (crosser_007_out_valid),             //          .valid
		.sink1_channel       (crosser_007_out_channel),           //          .channel
		.sink1_data          (crosser_007_out_data),              //          .data
		.sink1_startofpacket (crosser_007_out_startofpacket),     //          .startofpacket
		.sink1_endofpacket   (crosser_007_out_endofpacket)        //          .endofpacket
	);

	nios2VGA_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (crosser_008_out_ready),                 //     sink1.ready
		.sink1_valid          (crosser_008_out_valid),                 //          .valid
		.sink1_channel        (crosser_008_out_channel),               //          .channel
		.sink1_data           (crosser_008_out_data),                  //          .data
		.sink1_startofpacket  (crosser_008_out_startofpacket),         //          .startofpacket
		.sink1_endofpacket    (crosser_008_out_endofpacket),           //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (crosser_002_out_ready),                 //     sink6.ready
		.sink6_valid          (crosser_002_out_valid),                 //          .valid
		.sink6_channel        (crosser_002_out_channel),               //          .channel
		.sink6_data           (crosser_002_out_data),                  //          .data
		.sink6_startofpacket  (crosser_002_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket    (crosser_002_out_endofpacket),           //          .endofpacket
		.sink7_ready          (crosser_009_out_ready),                 //     sink7.ready
		.sink7_valid          (crosser_009_out_valid),                 //          .valid
		.sink7_channel        (crosser_009_out_channel),               //          .channel
		.sink7_data           (crosser_009_out_data),                  //          .data
		.sink7_startofpacket  (crosser_009_out_startofpacket),         //          .startofpacket
		.sink7_endofpacket    (crosser_009_out_endofpacket),           //          .endofpacket
		.sink8_ready          (crosser_003_out_ready),                 //     sink8.ready
		.sink8_valid          (crosser_003_out_valid),                 //          .valid
		.sink8_channel        (crosser_003_out_channel),               //          .channel
		.sink8_data           (crosser_003_out_data),                  //          .data
		.sink8_startofpacket  (crosser_003_out_startofpacket),         //          .startofpacket
		.sink8_endofpacket    (crosser_003_out_endofpacket),           //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (21),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk_clk),                           //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src1_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (21),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_001_src_data),            //          .data
		.out_channel          (width_adapter_001_src_channel),         //          .channel
		.out_valid            (width_adapter_001_src_valid),           //          .valid
		.out_ready            (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (81),
		.OUT_PKT_RESPONSE_STATUS_L     (80),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (21),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src7_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src7_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src7_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src7_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src7_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src7_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (21),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_003 (
		.clk                  (external_clocks_sys_clk_clk),           //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src0_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_003_src_data),            //          .data
		.out_channel          (width_adapter_003_src_channel),         //          .channel
		.out_valid            (width_adapter_003_src_valid),           //          .valid
		.out_ready            (width_adapter_003_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (21),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_004 (
		.clk                  (external_clocks_sys_clk_clk),           //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src2_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src2_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src2_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src2_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_004_src_data),            //          .data
		.out_channel          (width_adapter_004_src_channel),         //          .channel
		.out_valid            (width_adapter_004_src_valid),           //          .valid
		.out_ready            (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (81),
		.IN_PKT_RESPONSE_STATUS_L      (80),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (21),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_005 (
		.clk                  (external_clocks_sys_clk_clk),           //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_007_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_007_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_007_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_007_src0_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (external_clocks_sys_clk_clk),           //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src6_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (external_clocks_sys_clk_clk),           //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src8_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src8_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src8_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src8_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src8_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src8_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (external_clocks_sys_clk_clk),           //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (external_clocks_sys_clk_clk),           //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (91),
		.BITS_PER_SYMBOL     (91),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (external_clocks_sys_clk_clk),        //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset), // out_clk_reset.reset
		.in_ready          (width_adapter_src_ready),            //            in.ready
		.in_valid          (width_adapter_src_valid),            //              .valid
		.in_startofpacket  (width_adapter_src_startofpacket),    //              .startofpacket
		.in_endofpacket    (width_adapter_src_endofpacket),      //              .endofpacket
		.in_channel        (width_adapter_src_channel),          //              .channel
		.in_data           (width_adapter_src_data),             //              .data
		.out_ready         (crosser_004_out_ready),              //           out.ready
		.out_valid         (crosser_004_out_valid),              //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_004_out_channel),            //              .channel
		.out_data          (crosser_004_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (91),
		.BITS_PER_SYMBOL     (91),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (clk_clk),                             //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),      //  in_clk_reset.reset
		.out_clk           (external_clocks_sys_clk_clk),         //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),  // out_clk_reset.reset
		.in_ready          (width_adapter_001_src_ready),         //            in.ready
		.in_valid          (width_adapter_001_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_001_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_001_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_001_src_channel),       //              .channel
		.in_data           (width_adapter_001_src_data),          //              .data
		.out_ready         (crosser_005_out_ready),               //           out.ready
		.out_valid         (crosser_005_out_valid),               //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_005_out_channel),             //              .channel
		.out_data          (crosser_005_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (82),
		.BITS_PER_SYMBOL     (82),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (clk_clk),                             //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),      //  in_clk_reset.reset
		.out_clk           (external_clocks_sys_clk_clk),         //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),  // out_clk_reset.reset
		.in_ready          (width_adapter_002_src_ready),         //            in.ready
		.in_valid          (width_adapter_002_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_002_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_002_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_002_src_channel),       //              .channel
		.in_data           (width_adapter_002_src_data),          //              .data
		.out_ready         (crosser_006_out_ready),               //           out.ready
		.out_valid         (crosser_006_out_valid),               //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_006_out_channel),             //              .channel
		.out_data          (crosser_006_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (external_clocks_sys_clk_clk),         //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),  //  in_clk_reset.reset
		.out_clk           (clk_clk),                             //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),      // out_clk_reset.reset
		.in_ready          (width_adapter_003_src_ready),         //            in.ready
		.in_valid          (width_adapter_003_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_003_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_003_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_003_src_channel),       //              .channel
		.in_data           (width_adapter_003_src_data),          //              .data
		.out_ready         (crosser_007_out_ready),               //           out.ready
		.out_valid         (crosser_007_out_valid),               //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_007_out_channel),             //              .channel
		.out_data          (crosser_007_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_008 (
		.in_clk            (external_clocks_sys_clk_clk),         //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),  //  in_clk_reset.reset
		.out_clk           (clk_clk),                             //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),      // out_clk_reset.reset
		.in_ready          (width_adapter_004_src_ready),         //            in.ready
		.in_valid          (width_adapter_004_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_004_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_004_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_004_src_channel),       //              .channel
		.in_data           (width_adapter_004_src_data),          //              .data
		.out_ready         (crosser_008_out_ready),               //           out.ready
		.out_valid         (crosser_008_out_valid),               //              .valid
		.out_startofpacket (crosser_008_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_008_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_008_out_channel),             //              .channel
		.out_data          (crosser_008_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (21),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_009 (
		.in_clk            (external_clocks_sys_clk_clk),         //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),  //  in_clk_reset.reset
		.out_clk           (clk_clk),                             //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),      // out_clk_reset.reset
		.in_ready          (width_adapter_005_src_ready),         //            in.ready
		.in_valid          (width_adapter_005_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_005_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_005_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_005_src_channel),       //              .channel
		.in_data           (width_adapter_005_src_data),          //              .data
		.out_ready         (crosser_009_out_ready),               //           out.ready
		.out_valid         (crosser_009_out_valid),               //              .valid
		.out_startofpacket (crosser_009_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_009_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_009_out_channel),             //              .channel
		.out_data          (crosser_009_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	nios2VGA_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

endmodule
