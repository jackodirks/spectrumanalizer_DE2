library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

ENTITY fft_tld IS
PORT (
	adc_samples : IN STD_LOGIC_VECTOR(20479 DOWNTO 0);
	fft_samples : OUT STD_LOGIC_VECTOR(159 DOWNTO 0);
	samples_ready : IN STD_LOGIC := '0';	-- sampler has 2048 samples ready
	clk : IN STD_LOGIC := '0';
	fft_finished : OUT STD_LOGIC := '0';	-- the system is idle / can receive data
	busy : IN STD_LOGIC := '0';	-- receiving side status
	data_ready : OUT STD_LOGIC := '0' -- the FFT has data ready for output / cycle data
	);
END ENTITY;

ARCHITECTURE fft_tld OF fft_tld IS
	COMPONENT fft_peripheral IS
	PORT(
			X0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X16 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X17 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X18 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X19 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X20 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X21 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X22 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X23 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X24 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X25 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X26 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X27 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X28 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X29 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X30 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X31 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X32 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X33 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X34 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X35 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X36 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X37 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X38 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X39 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X40 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X41 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X42 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X43 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X44 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X45 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X46 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X47 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X48 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X49 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X50 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X51 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X52 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X53 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X54 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X55 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X56 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X57 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X58 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X59 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X60 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X61 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X62 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X63 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X64 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X65 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X66 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X67 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X68 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X69 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X70 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X71 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X72 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X73 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X74 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X75 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X76 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X77 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X78 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X79 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X80 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X81 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X82 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X83 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X84 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X85 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X86 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X87 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X88 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X89 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X90 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X91 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X92 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X93 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X94 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X95 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X96 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X97 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X98 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X99 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1048 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1049 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1050 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1051 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1052 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1053 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1054 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1055 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1056 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1057 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1058 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1059 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1060 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1061 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1062 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1063 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1064 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1065 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1066 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1067 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1068 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1069 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1070 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1071 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1072 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1073 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1074 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1075 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1076 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1077 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1078 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1079 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1080 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1081 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1082 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1083 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1084 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1085 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1086 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1087 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1088 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1089 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1090 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1091 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1092 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1093 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1094 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1095 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1096 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1097 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1098 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1099 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X1999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
			X2047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";	
		samples_ready : IN STD_LOGIC := '0';	-- sampler has 2048 samples ready
		clk : IN STD_LOGIC := '0';
		fft_finished : OUT STD_LOGIC := '0';	-- the system is idle / can receive data
	
		busy : IN STD_LOGIC := '0';	-- receiving side status
		data_ready : OUT STD_LOGIC := '0'; -- the FFT has data ready for output / cycle data
		
		-- data ouput for interfacing device 64 sets of 16 
		V0 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V1 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V2 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V3 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V4 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V5 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V6 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V7 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V8 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V9 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V10 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V11 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V12 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V13 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V14 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		V15 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000"
);
END COMPONENT;

BEGIN	

fft_peripheral_imp : fft_peripheral PORT MAP (
		X0 => adc_samples(9 DOWNTO 0),
	X1 => adc_samples(19 DOWNTO 10),
	X2 => adc_samples(29 DOWNTO 20),
	X3 => adc_samples(39 DOWNTO 30),
	X4 => adc_samples(49 DOWNTO 40),
	X5 => adc_samples(59 DOWNTO 50),
	X6 => adc_samples(69 DOWNTO 60),
	X7 => adc_samples(79 DOWNTO 70),
	X8 => adc_samples(89 DOWNTO 80),
	X9 => adc_samples(99 DOWNTO 90),
	X10 => adc_samples(109 DOWNTO 100),
	X11 => adc_samples(119 DOWNTO 110),
	X12 => adc_samples(129 DOWNTO 120),
	X13 => adc_samples(139 DOWNTO 130),
	X14 => adc_samples(149 DOWNTO 140),
	X15 => adc_samples(159 DOWNTO 150),
	X16 => adc_samples(169 DOWNTO 160),
	X17 => adc_samples(179 DOWNTO 170),
	X18 => adc_samples(189 DOWNTO 180),
	X19 => adc_samples(199 DOWNTO 190),
	X20 => adc_samples(209 DOWNTO 200),
	X21 => adc_samples(219 DOWNTO 210),
	X22 => adc_samples(229 DOWNTO 220),
	X23 => adc_samples(239 DOWNTO 230),
	X24 => adc_samples(249 DOWNTO 240),
	X25 => adc_samples(259 DOWNTO 250),
	X26 => adc_samples(269 DOWNTO 260),
	X27 => adc_samples(279 DOWNTO 270),
	X28 => adc_samples(289 DOWNTO 280),
	X29 => adc_samples(299 DOWNTO 290),
	X30 => adc_samples(309 DOWNTO 300),
	X31 => adc_samples(319 DOWNTO 310),
	X32 => adc_samples(329 DOWNTO 320),
	X33 => adc_samples(339 DOWNTO 330),
	X34 => adc_samples(349 DOWNTO 340),
	X35 => adc_samples(359 DOWNTO 350),
	X36 => adc_samples(369 DOWNTO 360),
	X37 => adc_samples(379 DOWNTO 370),
	X38 => adc_samples(389 DOWNTO 380),
	X39 => adc_samples(399 DOWNTO 390),
	X40 => adc_samples(409 DOWNTO 400),
	X41 => adc_samples(419 DOWNTO 410),
	X42 => adc_samples(429 DOWNTO 420),
	X43 => adc_samples(439 DOWNTO 430),
	X44 => adc_samples(449 DOWNTO 440),
	X45 => adc_samples(459 DOWNTO 450),
	X46 => adc_samples(469 DOWNTO 460),
	X47 => adc_samples(479 DOWNTO 470),
	X48 => adc_samples(489 DOWNTO 480),
	X49 => adc_samples(499 DOWNTO 490),
	X50 => adc_samples(509 DOWNTO 500),
	X51 => adc_samples(519 DOWNTO 510),
	X52 => adc_samples(529 DOWNTO 520),
	X53 => adc_samples(539 DOWNTO 530),
	X54 => adc_samples(549 DOWNTO 540),
	X55 => adc_samples(559 DOWNTO 550),
	X56 => adc_samples(569 DOWNTO 560),
	X57 => adc_samples(579 DOWNTO 570),
	X58 => adc_samples(589 DOWNTO 580),
	X59 => adc_samples(599 DOWNTO 590),
	X60 => adc_samples(609 DOWNTO 600),
	X61 => adc_samples(619 DOWNTO 610),
	X62 => adc_samples(629 DOWNTO 620),
	X63 => adc_samples(639 DOWNTO 630),
	X64 => adc_samples(649 DOWNTO 640),
	X65 => adc_samples(659 DOWNTO 650),
	X66 => adc_samples(669 DOWNTO 660),
	X67 => adc_samples(679 DOWNTO 670),
	X68 => adc_samples(689 DOWNTO 680),
	X69 => adc_samples(699 DOWNTO 690),
	X70 => adc_samples(709 DOWNTO 700),
	X71 => adc_samples(719 DOWNTO 710),
	X72 => adc_samples(729 DOWNTO 720),
	X73 => adc_samples(739 DOWNTO 730),
	X74 => adc_samples(749 DOWNTO 740),
	X75 => adc_samples(759 DOWNTO 750),
	X76 => adc_samples(769 DOWNTO 760),
	X77 => adc_samples(779 DOWNTO 770),
	X78 => adc_samples(789 DOWNTO 780),
	X79 => adc_samples(799 DOWNTO 790),
	X80 => adc_samples(809 DOWNTO 800),
	X81 => adc_samples(819 DOWNTO 810),
	X82 => adc_samples(829 DOWNTO 820),
	X83 => adc_samples(839 DOWNTO 830),
	X84 => adc_samples(849 DOWNTO 840),
	X85 => adc_samples(859 DOWNTO 850),
	X86 => adc_samples(869 DOWNTO 860),
	X87 => adc_samples(879 DOWNTO 870),
	X88 => adc_samples(889 DOWNTO 880),
	X89 => adc_samples(899 DOWNTO 890),
	X90 => adc_samples(909 DOWNTO 900),
	X91 => adc_samples(919 DOWNTO 910),
	X92 => adc_samples(929 DOWNTO 920),
	X93 => adc_samples(939 DOWNTO 930),
	X94 => adc_samples(949 DOWNTO 940),
	X95 => adc_samples(959 DOWNTO 950),
	X96 => adc_samples(969 DOWNTO 960),
	X97 => adc_samples(979 DOWNTO 970),
	X98 => adc_samples(989 DOWNTO 980),
	X99 => adc_samples(999 DOWNTO 990),
	X100 => adc_samples(1009 DOWNTO 1000),
	X101 => adc_samples(1019 DOWNTO 1010),
	X102 => adc_samples(1029 DOWNTO 1020),
	X103 => adc_samples(1039 DOWNTO 1030),
	X104 => adc_samples(1049 DOWNTO 1040),
	X105 => adc_samples(1059 DOWNTO 1050),
	X106 => adc_samples(1069 DOWNTO 1060),
	X107 => adc_samples(1079 DOWNTO 1070),
	X108 => adc_samples(1089 DOWNTO 1080),
	X109 => adc_samples(1099 DOWNTO 1090),
	X110 => adc_samples(1109 DOWNTO 1100),
	X111 => adc_samples(1119 DOWNTO 1110),
	X112 => adc_samples(1129 DOWNTO 1120),
	X113 => adc_samples(1139 DOWNTO 1130),
	X114 => adc_samples(1149 DOWNTO 1140),
	X115 => adc_samples(1159 DOWNTO 1150),
	X116 => adc_samples(1169 DOWNTO 1160),
	X117 => adc_samples(1179 DOWNTO 1170),
	X118 => adc_samples(1189 DOWNTO 1180),
	X119 => adc_samples(1199 DOWNTO 1190),
	X120 => adc_samples(1209 DOWNTO 1200),
	X121 => adc_samples(1219 DOWNTO 1210),
	X122 => adc_samples(1229 DOWNTO 1220),
	X123 => adc_samples(1239 DOWNTO 1230),
	X124 => adc_samples(1249 DOWNTO 1240),
	X125 => adc_samples(1259 DOWNTO 1250),
	X126 => adc_samples(1269 DOWNTO 1260),
	X127 => adc_samples(1279 DOWNTO 1270),
	X128 => adc_samples(1289 DOWNTO 1280),
	X129 => adc_samples(1299 DOWNTO 1290),
	X130 => adc_samples(1309 DOWNTO 1300),
	X131 => adc_samples(1319 DOWNTO 1310),
	X132 => adc_samples(1329 DOWNTO 1320),
	X133 => adc_samples(1339 DOWNTO 1330),
	X134 => adc_samples(1349 DOWNTO 1340),
	X135 => adc_samples(1359 DOWNTO 1350),
	X136 => adc_samples(1369 DOWNTO 1360),
	X137 => adc_samples(1379 DOWNTO 1370),
	X138 => adc_samples(1389 DOWNTO 1380),
	X139 => adc_samples(1399 DOWNTO 1390),
	X140 => adc_samples(1409 DOWNTO 1400),
	X141 => adc_samples(1419 DOWNTO 1410),
	X142 => adc_samples(1429 DOWNTO 1420),
	X143 => adc_samples(1439 DOWNTO 1430),
	X144 => adc_samples(1449 DOWNTO 1440),
	X145 => adc_samples(1459 DOWNTO 1450),
	X146 => adc_samples(1469 DOWNTO 1460),
	X147 => adc_samples(1479 DOWNTO 1470),
	X148 => adc_samples(1489 DOWNTO 1480),
	X149 => adc_samples(1499 DOWNTO 1490),
	X150 => adc_samples(1509 DOWNTO 1500),
	X151 => adc_samples(1519 DOWNTO 1510),
	X152 => adc_samples(1529 DOWNTO 1520),
	X153 => adc_samples(1539 DOWNTO 1530),
	X154 => adc_samples(1549 DOWNTO 1540),
	X155 => adc_samples(1559 DOWNTO 1550),
	X156 => adc_samples(1569 DOWNTO 1560),
	X157 => adc_samples(1579 DOWNTO 1570),
	X158 => adc_samples(1589 DOWNTO 1580),
	X159 => adc_samples(1599 DOWNTO 1590),
	X160 => adc_samples(1609 DOWNTO 1600),
	X161 => adc_samples(1619 DOWNTO 1610),
	X162 => adc_samples(1629 DOWNTO 1620),
	X163 => adc_samples(1639 DOWNTO 1630),
	X164 => adc_samples(1649 DOWNTO 1640),
	X165 => adc_samples(1659 DOWNTO 1650),
	X166 => adc_samples(1669 DOWNTO 1660),
	X167 => adc_samples(1679 DOWNTO 1670),
	X168 => adc_samples(1689 DOWNTO 1680),
	X169 => adc_samples(1699 DOWNTO 1690),
	X170 => adc_samples(1709 DOWNTO 1700),
	X171 => adc_samples(1719 DOWNTO 1710),
	X172 => adc_samples(1729 DOWNTO 1720),
	X173 => adc_samples(1739 DOWNTO 1730),
	X174 => adc_samples(1749 DOWNTO 1740),
	X175 => adc_samples(1759 DOWNTO 1750),
	X176 => adc_samples(1769 DOWNTO 1760),
	X177 => adc_samples(1779 DOWNTO 1770),
	X178 => adc_samples(1789 DOWNTO 1780),
	X179 => adc_samples(1799 DOWNTO 1790),
	X180 => adc_samples(1809 DOWNTO 1800),
	X181 => adc_samples(1819 DOWNTO 1810),
	X182 => adc_samples(1829 DOWNTO 1820),
	X183 => adc_samples(1839 DOWNTO 1830),
	X184 => adc_samples(1849 DOWNTO 1840),
	X185 => adc_samples(1859 DOWNTO 1850),
	X186 => adc_samples(1869 DOWNTO 1860),
	X187 => adc_samples(1879 DOWNTO 1870),
	X188 => adc_samples(1889 DOWNTO 1880),
	X189 => adc_samples(1899 DOWNTO 1890),
	X190 => adc_samples(1909 DOWNTO 1900),
	X191 => adc_samples(1919 DOWNTO 1910),
	X192 => adc_samples(1929 DOWNTO 1920),
	X193 => adc_samples(1939 DOWNTO 1930),
	X194 => adc_samples(1949 DOWNTO 1940),
	X195 => adc_samples(1959 DOWNTO 1950),
	X196 => adc_samples(1969 DOWNTO 1960),
	X197 => adc_samples(1979 DOWNTO 1970),
	X198 => adc_samples(1989 DOWNTO 1980),
	X199 => adc_samples(1999 DOWNTO 1990),
	X200 => adc_samples(2009 DOWNTO 2000),
	X201 => adc_samples(2019 DOWNTO 2010),
	X202 => adc_samples(2029 DOWNTO 2020),
	X203 => adc_samples(2039 DOWNTO 2030),
	X204 => adc_samples(2049 DOWNTO 2040),
	X205 => adc_samples(2059 DOWNTO 2050),
	X206 => adc_samples(2069 DOWNTO 2060),
	X207 => adc_samples(2079 DOWNTO 2070),
	X208 => adc_samples(2089 DOWNTO 2080),
	X209 => adc_samples(2099 DOWNTO 2090),
	X210 => adc_samples(2109 DOWNTO 2100),
	X211 => adc_samples(2119 DOWNTO 2110),
	X212 => adc_samples(2129 DOWNTO 2120),
	X213 => adc_samples(2139 DOWNTO 2130),
	X214 => adc_samples(2149 DOWNTO 2140),
	X215 => adc_samples(2159 DOWNTO 2150),
	X216 => adc_samples(2169 DOWNTO 2160),
	X217 => adc_samples(2179 DOWNTO 2170),
	X218 => adc_samples(2189 DOWNTO 2180),
	X219 => adc_samples(2199 DOWNTO 2190),
	X220 => adc_samples(2209 DOWNTO 2200),
	X221 => adc_samples(2219 DOWNTO 2210),
	X222 => adc_samples(2229 DOWNTO 2220),
	X223 => adc_samples(2239 DOWNTO 2230),
	X224 => adc_samples(2249 DOWNTO 2240),
	X225 => adc_samples(2259 DOWNTO 2250),
	X226 => adc_samples(2269 DOWNTO 2260),
	X227 => adc_samples(2279 DOWNTO 2270),
	X228 => adc_samples(2289 DOWNTO 2280),
	X229 => adc_samples(2299 DOWNTO 2290),
	X230 => adc_samples(2309 DOWNTO 2300),
	X231 => adc_samples(2319 DOWNTO 2310),
	X232 => adc_samples(2329 DOWNTO 2320),
	X233 => adc_samples(2339 DOWNTO 2330),
	X234 => adc_samples(2349 DOWNTO 2340),
	X235 => adc_samples(2359 DOWNTO 2350),
	X236 => adc_samples(2369 DOWNTO 2360),
	X237 => adc_samples(2379 DOWNTO 2370),
	X238 => adc_samples(2389 DOWNTO 2380),
	X239 => adc_samples(2399 DOWNTO 2390),
	X240 => adc_samples(2409 DOWNTO 2400),
	X241 => adc_samples(2419 DOWNTO 2410),
	X242 => adc_samples(2429 DOWNTO 2420),
	X243 => adc_samples(2439 DOWNTO 2430),
	X244 => adc_samples(2449 DOWNTO 2440),
	X245 => adc_samples(2459 DOWNTO 2450),
	X246 => adc_samples(2469 DOWNTO 2460),
	X247 => adc_samples(2479 DOWNTO 2470),
	X248 => adc_samples(2489 DOWNTO 2480),
	X249 => adc_samples(2499 DOWNTO 2490),
	X250 => adc_samples(2509 DOWNTO 2500),
	X251 => adc_samples(2519 DOWNTO 2510),
	X252 => adc_samples(2529 DOWNTO 2520),
	X253 => adc_samples(2539 DOWNTO 2530),
	X254 => adc_samples(2549 DOWNTO 2540),
	X255 => adc_samples(2559 DOWNTO 2550),
	X256 => adc_samples(2569 DOWNTO 2560),
	X257 => adc_samples(2579 DOWNTO 2570),
	X258 => adc_samples(2589 DOWNTO 2580),
	X259 => adc_samples(2599 DOWNTO 2590),
	X260 => adc_samples(2609 DOWNTO 2600),
	X261 => adc_samples(2619 DOWNTO 2610),
	X262 => adc_samples(2629 DOWNTO 2620),
	X263 => adc_samples(2639 DOWNTO 2630),
	X264 => adc_samples(2649 DOWNTO 2640),
	X265 => adc_samples(2659 DOWNTO 2650),
	X266 => adc_samples(2669 DOWNTO 2660),
	X267 => adc_samples(2679 DOWNTO 2670),
	X268 => adc_samples(2689 DOWNTO 2680),
	X269 => adc_samples(2699 DOWNTO 2690),
	X270 => adc_samples(2709 DOWNTO 2700),
	X271 => adc_samples(2719 DOWNTO 2710),
	X272 => adc_samples(2729 DOWNTO 2720),
	X273 => adc_samples(2739 DOWNTO 2730),
	X274 => adc_samples(2749 DOWNTO 2740),
	X275 => adc_samples(2759 DOWNTO 2750),
	X276 => adc_samples(2769 DOWNTO 2760),
	X277 => adc_samples(2779 DOWNTO 2770),
	X278 => adc_samples(2789 DOWNTO 2780),
	X279 => adc_samples(2799 DOWNTO 2790),
	X280 => adc_samples(2809 DOWNTO 2800),
	X281 => adc_samples(2819 DOWNTO 2810),
	X282 => adc_samples(2829 DOWNTO 2820),
	X283 => adc_samples(2839 DOWNTO 2830),
	X284 => adc_samples(2849 DOWNTO 2840),
	X285 => adc_samples(2859 DOWNTO 2850),
	X286 => adc_samples(2869 DOWNTO 2860),
	X287 => adc_samples(2879 DOWNTO 2870),
	X288 => adc_samples(2889 DOWNTO 2880),
	X289 => adc_samples(2899 DOWNTO 2890),
	X290 => adc_samples(2909 DOWNTO 2900),
	X291 => adc_samples(2919 DOWNTO 2910),
	X292 => adc_samples(2929 DOWNTO 2920),
	X293 => adc_samples(2939 DOWNTO 2930),
	X294 => adc_samples(2949 DOWNTO 2940),
	X295 => adc_samples(2959 DOWNTO 2950),
	X296 => adc_samples(2969 DOWNTO 2960),
	X297 => adc_samples(2979 DOWNTO 2970),
	X298 => adc_samples(2989 DOWNTO 2980),
	X299 => adc_samples(2999 DOWNTO 2990),
	X300 => adc_samples(3009 DOWNTO 3000),
	X301 => adc_samples(3019 DOWNTO 3010),
	X302 => adc_samples(3029 DOWNTO 3020),
	X303 => adc_samples(3039 DOWNTO 3030),
	X304 => adc_samples(3049 DOWNTO 3040),
	X305 => adc_samples(3059 DOWNTO 3050),
	X306 => adc_samples(3069 DOWNTO 3060),
	X307 => adc_samples(3079 DOWNTO 3070),
	X308 => adc_samples(3089 DOWNTO 3080),
	X309 => adc_samples(3099 DOWNTO 3090),
	X310 => adc_samples(3109 DOWNTO 3100),
	X311 => adc_samples(3119 DOWNTO 3110),
	X312 => adc_samples(3129 DOWNTO 3120),
	X313 => adc_samples(3139 DOWNTO 3130),
	X314 => adc_samples(3149 DOWNTO 3140),
	X315 => adc_samples(3159 DOWNTO 3150),
	X316 => adc_samples(3169 DOWNTO 3160),
	X317 => adc_samples(3179 DOWNTO 3170),
	X318 => adc_samples(3189 DOWNTO 3180),
	X319 => adc_samples(3199 DOWNTO 3190),
	X320 => adc_samples(3209 DOWNTO 3200),
	X321 => adc_samples(3219 DOWNTO 3210),
	X322 => adc_samples(3229 DOWNTO 3220),
	X323 => adc_samples(3239 DOWNTO 3230),
	X324 => adc_samples(3249 DOWNTO 3240),
	X325 => adc_samples(3259 DOWNTO 3250),
	X326 => adc_samples(3269 DOWNTO 3260),
	X327 => adc_samples(3279 DOWNTO 3270),
	X328 => adc_samples(3289 DOWNTO 3280),
	X329 => adc_samples(3299 DOWNTO 3290),
	X330 => adc_samples(3309 DOWNTO 3300),
	X331 => adc_samples(3319 DOWNTO 3310),
	X332 => adc_samples(3329 DOWNTO 3320),
	X333 => adc_samples(3339 DOWNTO 3330),
	X334 => adc_samples(3349 DOWNTO 3340),
	X335 => adc_samples(3359 DOWNTO 3350),
	X336 => adc_samples(3369 DOWNTO 3360),
	X337 => adc_samples(3379 DOWNTO 3370),
	X338 => adc_samples(3389 DOWNTO 3380),
	X339 => adc_samples(3399 DOWNTO 3390),
	X340 => adc_samples(3409 DOWNTO 3400),
	X341 => adc_samples(3419 DOWNTO 3410),
	X342 => adc_samples(3429 DOWNTO 3420),
	X343 => adc_samples(3439 DOWNTO 3430),
	X344 => adc_samples(3449 DOWNTO 3440),
	X345 => adc_samples(3459 DOWNTO 3450),
	X346 => adc_samples(3469 DOWNTO 3460),
	X347 => adc_samples(3479 DOWNTO 3470),
	X348 => adc_samples(3489 DOWNTO 3480),
	X349 => adc_samples(3499 DOWNTO 3490),
	X350 => adc_samples(3509 DOWNTO 3500),
	X351 => adc_samples(3519 DOWNTO 3510),
	X352 => adc_samples(3529 DOWNTO 3520),
	X353 => adc_samples(3539 DOWNTO 3530),
	X354 => adc_samples(3549 DOWNTO 3540),
	X355 => adc_samples(3559 DOWNTO 3550),
	X356 => adc_samples(3569 DOWNTO 3560),
	X357 => adc_samples(3579 DOWNTO 3570),
	X358 => adc_samples(3589 DOWNTO 3580),
	X359 => adc_samples(3599 DOWNTO 3590),
	X360 => adc_samples(3609 DOWNTO 3600),
	X361 => adc_samples(3619 DOWNTO 3610),
	X362 => adc_samples(3629 DOWNTO 3620),
	X363 => adc_samples(3639 DOWNTO 3630),
	X364 => adc_samples(3649 DOWNTO 3640),
	X365 => adc_samples(3659 DOWNTO 3650),
	X366 => adc_samples(3669 DOWNTO 3660),
	X367 => adc_samples(3679 DOWNTO 3670),
	X368 => adc_samples(3689 DOWNTO 3680),
	X369 => adc_samples(3699 DOWNTO 3690),
	X370 => adc_samples(3709 DOWNTO 3700),
	X371 => adc_samples(3719 DOWNTO 3710),
	X372 => adc_samples(3729 DOWNTO 3720),
	X373 => adc_samples(3739 DOWNTO 3730),
	X374 => adc_samples(3749 DOWNTO 3740),
	X375 => adc_samples(3759 DOWNTO 3750),
	X376 => adc_samples(3769 DOWNTO 3760),
	X377 => adc_samples(3779 DOWNTO 3770),
	X378 => adc_samples(3789 DOWNTO 3780),
	X379 => adc_samples(3799 DOWNTO 3790),
	X380 => adc_samples(3809 DOWNTO 3800),
	X381 => adc_samples(3819 DOWNTO 3810),
	X382 => adc_samples(3829 DOWNTO 3820),
	X383 => adc_samples(3839 DOWNTO 3830),
	X384 => adc_samples(3849 DOWNTO 3840),
	X385 => adc_samples(3859 DOWNTO 3850),
	X386 => adc_samples(3869 DOWNTO 3860),
	X387 => adc_samples(3879 DOWNTO 3870),
	X388 => adc_samples(3889 DOWNTO 3880),
	X389 => adc_samples(3899 DOWNTO 3890),
	X390 => adc_samples(3909 DOWNTO 3900),
	X391 => adc_samples(3919 DOWNTO 3910),
	X392 => adc_samples(3929 DOWNTO 3920),
	X393 => adc_samples(3939 DOWNTO 3930),
	X394 => adc_samples(3949 DOWNTO 3940),
	X395 => adc_samples(3959 DOWNTO 3950),
	X396 => adc_samples(3969 DOWNTO 3960),
	X397 => adc_samples(3979 DOWNTO 3970),
	X398 => adc_samples(3989 DOWNTO 3980),
	X399 => adc_samples(3999 DOWNTO 3990),
	X400 => adc_samples(4009 DOWNTO 4000),
	X401 => adc_samples(4019 DOWNTO 4010),
	X402 => adc_samples(4029 DOWNTO 4020),
	X403 => adc_samples(4039 DOWNTO 4030),
	X404 => adc_samples(4049 DOWNTO 4040),
	X405 => adc_samples(4059 DOWNTO 4050),
	X406 => adc_samples(4069 DOWNTO 4060),
	X407 => adc_samples(4079 DOWNTO 4070),
	X408 => adc_samples(4089 DOWNTO 4080),
	X409 => adc_samples(4099 DOWNTO 4090),
	X410 => adc_samples(4109 DOWNTO 4100),
	X411 => adc_samples(4119 DOWNTO 4110),
	X412 => adc_samples(4129 DOWNTO 4120),
	X413 => adc_samples(4139 DOWNTO 4130),
	X414 => adc_samples(4149 DOWNTO 4140),
	X415 => adc_samples(4159 DOWNTO 4150),
	X416 => adc_samples(4169 DOWNTO 4160),
	X417 => adc_samples(4179 DOWNTO 4170),
	X418 => adc_samples(4189 DOWNTO 4180),
	X419 => adc_samples(4199 DOWNTO 4190),
	X420 => adc_samples(4209 DOWNTO 4200),
	X421 => adc_samples(4219 DOWNTO 4210),
	X422 => adc_samples(4229 DOWNTO 4220),
	X423 => adc_samples(4239 DOWNTO 4230),
	X424 => adc_samples(4249 DOWNTO 4240),
	X425 => adc_samples(4259 DOWNTO 4250),
	X426 => adc_samples(4269 DOWNTO 4260),
	X427 => adc_samples(4279 DOWNTO 4270),
	X428 => adc_samples(4289 DOWNTO 4280),
	X429 => adc_samples(4299 DOWNTO 4290),
	X430 => adc_samples(4309 DOWNTO 4300),
	X431 => adc_samples(4319 DOWNTO 4310),
	X432 => adc_samples(4329 DOWNTO 4320),
	X433 => adc_samples(4339 DOWNTO 4330),
	X434 => adc_samples(4349 DOWNTO 4340),
	X435 => adc_samples(4359 DOWNTO 4350),
	X436 => adc_samples(4369 DOWNTO 4360),
	X437 => adc_samples(4379 DOWNTO 4370),
	X438 => adc_samples(4389 DOWNTO 4380),
	X439 => adc_samples(4399 DOWNTO 4390),
	X440 => adc_samples(4409 DOWNTO 4400),
	X441 => adc_samples(4419 DOWNTO 4410),
	X442 => adc_samples(4429 DOWNTO 4420),
	X443 => adc_samples(4439 DOWNTO 4430),
	X444 => adc_samples(4449 DOWNTO 4440),
	X445 => adc_samples(4459 DOWNTO 4450),
	X446 => adc_samples(4469 DOWNTO 4460),
	X447 => adc_samples(4479 DOWNTO 4470),
	X448 => adc_samples(4489 DOWNTO 4480),
	X449 => adc_samples(4499 DOWNTO 4490),
	X450 => adc_samples(4509 DOWNTO 4500),
	X451 => adc_samples(4519 DOWNTO 4510),
	X452 => adc_samples(4529 DOWNTO 4520),
	X453 => adc_samples(4539 DOWNTO 4530),
	X454 => adc_samples(4549 DOWNTO 4540),
	X455 => adc_samples(4559 DOWNTO 4550),
	X456 => adc_samples(4569 DOWNTO 4560),
	X457 => adc_samples(4579 DOWNTO 4570),
	X458 => adc_samples(4589 DOWNTO 4580),
	X459 => adc_samples(4599 DOWNTO 4590),
	X460 => adc_samples(4609 DOWNTO 4600),
	X461 => adc_samples(4619 DOWNTO 4610),
	X462 => adc_samples(4629 DOWNTO 4620),
	X463 => adc_samples(4639 DOWNTO 4630),
	X464 => adc_samples(4649 DOWNTO 4640),
	X465 => adc_samples(4659 DOWNTO 4650),
	X466 => adc_samples(4669 DOWNTO 4660),
	X467 => adc_samples(4679 DOWNTO 4670),
	X468 => adc_samples(4689 DOWNTO 4680),
	X469 => adc_samples(4699 DOWNTO 4690),
	X470 => adc_samples(4709 DOWNTO 4700),
	X471 => adc_samples(4719 DOWNTO 4710),
	X472 => adc_samples(4729 DOWNTO 4720),
	X473 => adc_samples(4739 DOWNTO 4730),
	X474 => adc_samples(4749 DOWNTO 4740),
	X475 => adc_samples(4759 DOWNTO 4750),
	X476 => adc_samples(4769 DOWNTO 4760),
	X477 => adc_samples(4779 DOWNTO 4770),
	X478 => adc_samples(4789 DOWNTO 4780),
	X479 => adc_samples(4799 DOWNTO 4790),
	X480 => adc_samples(4809 DOWNTO 4800),
	X481 => adc_samples(4819 DOWNTO 4810),
	X482 => adc_samples(4829 DOWNTO 4820),
	X483 => adc_samples(4839 DOWNTO 4830),
	X484 => adc_samples(4849 DOWNTO 4840),
	X485 => adc_samples(4859 DOWNTO 4850),
	X486 => adc_samples(4869 DOWNTO 4860),
	X487 => adc_samples(4879 DOWNTO 4870),
	X488 => adc_samples(4889 DOWNTO 4880),
	X489 => adc_samples(4899 DOWNTO 4890),
	X490 => adc_samples(4909 DOWNTO 4900),
	X491 => adc_samples(4919 DOWNTO 4910),
	X492 => adc_samples(4929 DOWNTO 4920),
	X493 => adc_samples(4939 DOWNTO 4930),
	X494 => adc_samples(4949 DOWNTO 4940),
	X495 => adc_samples(4959 DOWNTO 4950),
	X496 => adc_samples(4969 DOWNTO 4960),
	X497 => adc_samples(4979 DOWNTO 4970),
	X498 => adc_samples(4989 DOWNTO 4980),
	X499 => adc_samples(4999 DOWNTO 4990),
	X500 => adc_samples(5009 DOWNTO 5000),
	X501 => adc_samples(5019 DOWNTO 5010),
	X502 => adc_samples(5029 DOWNTO 5020),
	X503 => adc_samples(5039 DOWNTO 5030),
	X504 => adc_samples(5049 DOWNTO 5040),
	X505 => adc_samples(5059 DOWNTO 5050),
	X506 => adc_samples(5069 DOWNTO 5060),
	X507 => adc_samples(5079 DOWNTO 5070),
	X508 => adc_samples(5089 DOWNTO 5080),
	X509 => adc_samples(5099 DOWNTO 5090),
	X510 => adc_samples(5109 DOWNTO 5100),
	X511 => adc_samples(5119 DOWNTO 5110),
	X512 => adc_samples(5129 DOWNTO 5120),
	X513 => adc_samples(5139 DOWNTO 5130),
	X514 => adc_samples(5149 DOWNTO 5140),
	X515 => adc_samples(5159 DOWNTO 5150),
	X516 => adc_samples(5169 DOWNTO 5160),
	X517 => adc_samples(5179 DOWNTO 5170),
	X518 => adc_samples(5189 DOWNTO 5180),
	X519 => adc_samples(5199 DOWNTO 5190),
	X520 => adc_samples(5209 DOWNTO 5200),
	X521 => adc_samples(5219 DOWNTO 5210),
	X522 => adc_samples(5229 DOWNTO 5220),
	X523 => adc_samples(5239 DOWNTO 5230),
	X524 => adc_samples(5249 DOWNTO 5240),
	X525 => adc_samples(5259 DOWNTO 5250),
	X526 => adc_samples(5269 DOWNTO 5260),
	X527 => adc_samples(5279 DOWNTO 5270),
	X528 => adc_samples(5289 DOWNTO 5280),
	X529 => adc_samples(5299 DOWNTO 5290),
	X530 => adc_samples(5309 DOWNTO 5300),
	X531 => adc_samples(5319 DOWNTO 5310),
	X532 => adc_samples(5329 DOWNTO 5320),
	X533 => adc_samples(5339 DOWNTO 5330),
	X534 => adc_samples(5349 DOWNTO 5340),
	X535 => adc_samples(5359 DOWNTO 5350),
	X536 => adc_samples(5369 DOWNTO 5360),
	X537 => adc_samples(5379 DOWNTO 5370),
	X538 => adc_samples(5389 DOWNTO 5380),
	X539 => adc_samples(5399 DOWNTO 5390),
	X540 => adc_samples(5409 DOWNTO 5400),
	X541 => adc_samples(5419 DOWNTO 5410),
	X542 => adc_samples(5429 DOWNTO 5420),
	X543 => adc_samples(5439 DOWNTO 5430),
	X544 => adc_samples(5449 DOWNTO 5440),
	X545 => adc_samples(5459 DOWNTO 5450),
	X546 => adc_samples(5469 DOWNTO 5460),
	X547 => adc_samples(5479 DOWNTO 5470),
	X548 => adc_samples(5489 DOWNTO 5480),
	X549 => adc_samples(5499 DOWNTO 5490),
	X550 => adc_samples(5509 DOWNTO 5500),
	X551 => adc_samples(5519 DOWNTO 5510),
	X552 => adc_samples(5529 DOWNTO 5520),
	X553 => adc_samples(5539 DOWNTO 5530),
	X554 => adc_samples(5549 DOWNTO 5540),
	X555 => adc_samples(5559 DOWNTO 5550),
	X556 => adc_samples(5569 DOWNTO 5560),
	X557 => adc_samples(5579 DOWNTO 5570),
	X558 => adc_samples(5589 DOWNTO 5580),
	X559 => adc_samples(5599 DOWNTO 5590),
	X560 => adc_samples(5609 DOWNTO 5600),
	X561 => adc_samples(5619 DOWNTO 5610),
	X562 => adc_samples(5629 DOWNTO 5620),
	X563 => adc_samples(5639 DOWNTO 5630),
	X564 => adc_samples(5649 DOWNTO 5640),
	X565 => adc_samples(5659 DOWNTO 5650),
	X566 => adc_samples(5669 DOWNTO 5660),
	X567 => adc_samples(5679 DOWNTO 5670),
	X568 => adc_samples(5689 DOWNTO 5680),
	X569 => adc_samples(5699 DOWNTO 5690),
	X570 => adc_samples(5709 DOWNTO 5700),
	X571 => adc_samples(5719 DOWNTO 5710),
	X572 => adc_samples(5729 DOWNTO 5720),
	X573 => adc_samples(5739 DOWNTO 5730),
	X574 => adc_samples(5749 DOWNTO 5740),
	X575 => adc_samples(5759 DOWNTO 5750),
	X576 => adc_samples(5769 DOWNTO 5760),
	X577 => adc_samples(5779 DOWNTO 5770),
	X578 => adc_samples(5789 DOWNTO 5780),
	X579 => adc_samples(5799 DOWNTO 5790),
	X580 => adc_samples(5809 DOWNTO 5800),
	X581 => adc_samples(5819 DOWNTO 5810),
	X582 => adc_samples(5829 DOWNTO 5820),
	X583 => adc_samples(5839 DOWNTO 5830),
	X584 => adc_samples(5849 DOWNTO 5840),
	X585 => adc_samples(5859 DOWNTO 5850),
	X586 => adc_samples(5869 DOWNTO 5860),
	X587 => adc_samples(5879 DOWNTO 5870),
	X588 => adc_samples(5889 DOWNTO 5880),
	X589 => adc_samples(5899 DOWNTO 5890),
	X590 => adc_samples(5909 DOWNTO 5900),
	X591 => adc_samples(5919 DOWNTO 5910),
	X592 => adc_samples(5929 DOWNTO 5920),
	X593 => adc_samples(5939 DOWNTO 5930),
	X594 => adc_samples(5949 DOWNTO 5940),
	X595 => adc_samples(5959 DOWNTO 5950),
	X596 => adc_samples(5969 DOWNTO 5960),
	X597 => adc_samples(5979 DOWNTO 5970),
	X598 => adc_samples(5989 DOWNTO 5980),
	X599 => adc_samples(5999 DOWNTO 5990),
	X600 => adc_samples(6009 DOWNTO 6000),
	X601 => adc_samples(6019 DOWNTO 6010),
	X602 => adc_samples(6029 DOWNTO 6020),
	X603 => adc_samples(6039 DOWNTO 6030),
	X604 => adc_samples(6049 DOWNTO 6040),
	X605 => adc_samples(6059 DOWNTO 6050),
	X606 => adc_samples(6069 DOWNTO 6060),
	X607 => adc_samples(6079 DOWNTO 6070),
	X608 => adc_samples(6089 DOWNTO 6080),
	X609 => adc_samples(6099 DOWNTO 6090),
	X610 => adc_samples(6109 DOWNTO 6100),
	X611 => adc_samples(6119 DOWNTO 6110),
	X612 => adc_samples(6129 DOWNTO 6120),
	X613 => adc_samples(6139 DOWNTO 6130),
	X614 => adc_samples(6149 DOWNTO 6140),
	X615 => adc_samples(6159 DOWNTO 6150),
	X616 => adc_samples(6169 DOWNTO 6160),
	X617 => adc_samples(6179 DOWNTO 6170),
	X618 => adc_samples(6189 DOWNTO 6180),
	X619 => adc_samples(6199 DOWNTO 6190),
	X620 => adc_samples(6209 DOWNTO 6200),
	X621 => adc_samples(6219 DOWNTO 6210),
	X622 => adc_samples(6229 DOWNTO 6220),
	X623 => adc_samples(6239 DOWNTO 6230),
	X624 => adc_samples(6249 DOWNTO 6240),
	X625 => adc_samples(6259 DOWNTO 6250),
	X626 => adc_samples(6269 DOWNTO 6260),
	X627 => adc_samples(6279 DOWNTO 6270),
	X628 => adc_samples(6289 DOWNTO 6280),
	X629 => adc_samples(6299 DOWNTO 6290),
	X630 => adc_samples(6309 DOWNTO 6300),
	X631 => adc_samples(6319 DOWNTO 6310),
	X632 => adc_samples(6329 DOWNTO 6320),
	X633 => adc_samples(6339 DOWNTO 6330),
	X634 => adc_samples(6349 DOWNTO 6340),
	X635 => adc_samples(6359 DOWNTO 6350),
	X636 => adc_samples(6369 DOWNTO 6360),
	X637 => adc_samples(6379 DOWNTO 6370),
	X638 => adc_samples(6389 DOWNTO 6380),
	X639 => adc_samples(6399 DOWNTO 6390),
	X640 => adc_samples(6409 DOWNTO 6400),
	X641 => adc_samples(6419 DOWNTO 6410),
	X642 => adc_samples(6429 DOWNTO 6420),
	X643 => adc_samples(6439 DOWNTO 6430),
	X644 => adc_samples(6449 DOWNTO 6440),
	X645 => adc_samples(6459 DOWNTO 6450),
	X646 => adc_samples(6469 DOWNTO 6460),
	X647 => adc_samples(6479 DOWNTO 6470),
	X648 => adc_samples(6489 DOWNTO 6480),
	X649 => adc_samples(6499 DOWNTO 6490),
	X650 => adc_samples(6509 DOWNTO 6500),
	X651 => adc_samples(6519 DOWNTO 6510),
	X652 => adc_samples(6529 DOWNTO 6520),
	X653 => adc_samples(6539 DOWNTO 6530),
	X654 => adc_samples(6549 DOWNTO 6540),
	X655 => adc_samples(6559 DOWNTO 6550),
	X656 => adc_samples(6569 DOWNTO 6560),
	X657 => adc_samples(6579 DOWNTO 6570),
	X658 => adc_samples(6589 DOWNTO 6580),
	X659 => adc_samples(6599 DOWNTO 6590),
	X660 => adc_samples(6609 DOWNTO 6600),
	X661 => adc_samples(6619 DOWNTO 6610),
	X662 => adc_samples(6629 DOWNTO 6620),
	X663 => adc_samples(6639 DOWNTO 6630),
	X664 => adc_samples(6649 DOWNTO 6640),
	X665 => adc_samples(6659 DOWNTO 6650),
	X666 => adc_samples(6669 DOWNTO 6660),
	X667 => adc_samples(6679 DOWNTO 6670),
	X668 => adc_samples(6689 DOWNTO 6680),
	X669 => adc_samples(6699 DOWNTO 6690),
	X670 => adc_samples(6709 DOWNTO 6700),
	X671 => adc_samples(6719 DOWNTO 6710),
	X672 => adc_samples(6729 DOWNTO 6720),
	X673 => adc_samples(6739 DOWNTO 6730),
	X674 => adc_samples(6749 DOWNTO 6740),
	X675 => adc_samples(6759 DOWNTO 6750),
	X676 => adc_samples(6769 DOWNTO 6760),
	X677 => adc_samples(6779 DOWNTO 6770),
	X678 => adc_samples(6789 DOWNTO 6780),
	X679 => adc_samples(6799 DOWNTO 6790),
	X680 => adc_samples(6809 DOWNTO 6800),
	X681 => adc_samples(6819 DOWNTO 6810),
	X682 => adc_samples(6829 DOWNTO 6820),
	X683 => adc_samples(6839 DOWNTO 6830),
	X684 => adc_samples(6849 DOWNTO 6840),
	X685 => adc_samples(6859 DOWNTO 6850),
	X686 => adc_samples(6869 DOWNTO 6860),
	X687 => adc_samples(6879 DOWNTO 6870),
	X688 => adc_samples(6889 DOWNTO 6880),
	X689 => adc_samples(6899 DOWNTO 6890),
	X690 => adc_samples(6909 DOWNTO 6900),
	X691 => adc_samples(6919 DOWNTO 6910),
	X692 => adc_samples(6929 DOWNTO 6920),
	X693 => adc_samples(6939 DOWNTO 6930),
	X694 => adc_samples(6949 DOWNTO 6940),
	X695 => adc_samples(6959 DOWNTO 6950),
	X696 => adc_samples(6969 DOWNTO 6960),
	X697 => adc_samples(6979 DOWNTO 6970),
	X698 => adc_samples(6989 DOWNTO 6980),
	X699 => adc_samples(6999 DOWNTO 6990),
	X700 => adc_samples(7009 DOWNTO 7000),
	X701 => adc_samples(7019 DOWNTO 7010),
	X702 => adc_samples(7029 DOWNTO 7020),
	X703 => adc_samples(7039 DOWNTO 7030),
	X704 => adc_samples(7049 DOWNTO 7040),
	X705 => adc_samples(7059 DOWNTO 7050),
	X706 => adc_samples(7069 DOWNTO 7060),
	X707 => adc_samples(7079 DOWNTO 7070),
	X708 => adc_samples(7089 DOWNTO 7080),
	X709 => adc_samples(7099 DOWNTO 7090),
	X710 => adc_samples(7109 DOWNTO 7100),
	X711 => adc_samples(7119 DOWNTO 7110),
	X712 => adc_samples(7129 DOWNTO 7120),
	X713 => adc_samples(7139 DOWNTO 7130),
	X714 => adc_samples(7149 DOWNTO 7140),
	X715 => adc_samples(7159 DOWNTO 7150),
	X716 => adc_samples(7169 DOWNTO 7160),
	X717 => adc_samples(7179 DOWNTO 7170),
	X718 => adc_samples(7189 DOWNTO 7180),
	X719 => adc_samples(7199 DOWNTO 7190),
	X720 => adc_samples(7209 DOWNTO 7200),
	X721 => adc_samples(7219 DOWNTO 7210),
	X722 => adc_samples(7229 DOWNTO 7220),
	X723 => adc_samples(7239 DOWNTO 7230),
	X724 => adc_samples(7249 DOWNTO 7240),
	X725 => adc_samples(7259 DOWNTO 7250),
	X726 => adc_samples(7269 DOWNTO 7260),
	X727 => adc_samples(7279 DOWNTO 7270),
	X728 => adc_samples(7289 DOWNTO 7280),
	X729 => adc_samples(7299 DOWNTO 7290),
	X730 => adc_samples(7309 DOWNTO 7300),
	X731 => adc_samples(7319 DOWNTO 7310),
	X732 => adc_samples(7329 DOWNTO 7320),
	X733 => adc_samples(7339 DOWNTO 7330),
	X734 => adc_samples(7349 DOWNTO 7340),
	X735 => adc_samples(7359 DOWNTO 7350),
	X736 => adc_samples(7369 DOWNTO 7360),
	X737 => adc_samples(7379 DOWNTO 7370),
	X738 => adc_samples(7389 DOWNTO 7380),
	X739 => adc_samples(7399 DOWNTO 7390),
	X740 => adc_samples(7409 DOWNTO 7400),
	X741 => adc_samples(7419 DOWNTO 7410),
	X742 => adc_samples(7429 DOWNTO 7420),
	X743 => adc_samples(7439 DOWNTO 7430),
	X744 => adc_samples(7449 DOWNTO 7440),
	X745 => adc_samples(7459 DOWNTO 7450),
	X746 => adc_samples(7469 DOWNTO 7460),
	X747 => adc_samples(7479 DOWNTO 7470),
	X748 => adc_samples(7489 DOWNTO 7480),
	X749 => adc_samples(7499 DOWNTO 7490),
	X750 => adc_samples(7509 DOWNTO 7500),
	X751 => adc_samples(7519 DOWNTO 7510),
	X752 => adc_samples(7529 DOWNTO 7520),
	X753 => adc_samples(7539 DOWNTO 7530),
	X754 => adc_samples(7549 DOWNTO 7540),
	X755 => adc_samples(7559 DOWNTO 7550),
	X756 => adc_samples(7569 DOWNTO 7560),
	X757 => adc_samples(7579 DOWNTO 7570),
	X758 => adc_samples(7589 DOWNTO 7580),
	X759 => adc_samples(7599 DOWNTO 7590),
	X760 => adc_samples(7609 DOWNTO 7600),
	X761 => adc_samples(7619 DOWNTO 7610),
	X762 => adc_samples(7629 DOWNTO 7620),
	X763 => adc_samples(7639 DOWNTO 7630),
	X764 => adc_samples(7649 DOWNTO 7640),
	X765 => adc_samples(7659 DOWNTO 7650),
	X766 => adc_samples(7669 DOWNTO 7660),
	X767 => adc_samples(7679 DOWNTO 7670),
	X768 => adc_samples(7689 DOWNTO 7680),
	X769 => adc_samples(7699 DOWNTO 7690),
	X770 => adc_samples(7709 DOWNTO 7700),
	X771 => adc_samples(7719 DOWNTO 7710),
	X772 => adc_samples(7729 DOWNTO 7720),
	X773 => adc_samples(7739 DOWNTO 7730),
	X774 => adc_samples(7749 DOWNTO 7740),
	X775 => adc_samples(7759 DOWNTO 7750),
	X776 => adc_samples(7769 DOWNTO 7760),
	X777 => adc_samples(7779 DOWNTO 7770),
	X778 => adc_samples(7789 DOWNTO 7780),
	X779 => adc_samples(7799 DOWNTO 7790),
	X780 => adc_samples(7809 DOWNTO 7800),
	X781 => adc_samples(7819 DOWNTO 7810),
	X782 => adc_samples(7829 DOWNTO 7820),
	X783 => adc_samples(7839 DOWNTO 7830),
	X784 => adc_samples(7849 DOWNTO 7840),
	X785 => adc_samples(7859 DOWNTO 7850),
	X786 => adc_samples(7869 DOWNTO 7860),
	X787 => adc_samples(7879 DOWNTO 7870),
	X788 => adc_samples(7889 DOWNTO 7880),
	X789 => adc_samples(7899 DOWNTO 7890),
	X790 => adc_samples(7909 DOWNTO 7900),
	X791 => adc_samples(7919 DOWNTO 7910),
	X792 => adc_samples(7929 DOWNTO 7920),
	X793 => adc_samples(7939 DOWNTO 7930),
	X794 => adc_samples(7949 DOWNTO 7940),
	X795 => adc_samples(7959 DOWNTO 7950),
	X796 => adc_samples(7969 DOWNTO 7960),
	X797 => adc_samples(7979 DOWNTO 7970),
	X798 => adc_samples(7989 DOWNTO 7980),
	X799 => adc_samples(7999 DOWNTO 7990),
	X800 => adc_samples(8009 DOWNTO 8000),
	X801 => adc_samples(8019 DOWNTO 8010),
	X802 => adc_samples(8029 DOWNTO 8020),
	X803 => adc_samples(8039 DOWNTO 8030),
	X804 => adc_samples(8049 DOWNTO 8040),
	X805 => adc_samples(8059 DOWNTO 8050),
	X806 => adc_samples(8069 DOWNTO 8060),
	X807 => adc_samples(8079 DOWNTO 8070),
	X808 => adc_samples(8089 DOWNTO 8080),
	X809 => adc_samples(8099 DOWNTO 8090),
	X810 => adc_samples(8109 DOWNTO 8100),
	X811 => adc_samples(8119 DOWNTO 8110),
	X812 => adc_samples(8129 DOWNTO 8120),
	X813 => adc_samples(8139 DOWNTO 8130),
	X814 => adc_samples(8149 DOWNTO 8140),
	X815 => adc_samples(8159 DOWNTO 8150),
	X816 => adc_samples(8169 DOWNTO 8160),
	X817 => adc_samples(8179 DOWNTO 8170),
	X818 => adc_samples(8189 DOWNTO 8180),
	X819 => adc_samples(8199 DOWNTO 8190),
	X820 => adc_samples(8209 DOWNTO 8200),
	X821 => adc_samples(8219 DOWNTO 8210),
	X822 => adc_samples(8229 DOWNTO 8220),
	X823 => adc_samples(8239 DOWNTO 8230),
	X824 => adc_samples(8249 DOWNTO 8240),
	X825 => adc_samples(8259 DOWNTO 8250),
	X826 => adc_samples(8269 DOWNTO 8260),
	X827 => adc_samples(8279 DOWNTO 8270),
	X828 => adc_samples(8289 DOWNTO 8280),
	X829 => adc_samples(8299 DOWNTO 8290),
	X830 => adc_samples(8309 DOWNTO 8300),
	X831 => adc_samples(8319 DOWNTO 8310),
	X832 => adc_samples(8329 DOWNTO 8320),
	X833 => adc_samples(8339 DOWNTO 8330),
	X834 => adc_samples(8349 DOWNTO 8340),
	X835 => adc_samples(8359 DOWNTO 8350),
	X836 => adc_samples(8369 DOWNTO 8360),
	X837 => adc_samples(8379 DOWNTO 8370),
	X838 => adc_samples(8389 DOWNTO 8380),
	X839 => adc_samples(8399 DOWNTO 8390),
	X840 => adc_samples(8409 DOWNTO 8400),
	X841 => adc_samples(8419 DOWNTO 8410),
	X842 => adc_samples(8429 DOWNTO 8420),
	X843 => adc_samples(8439 DOWNTO 8430),
	X844 => adc_samples(8449 DOWNTO 8440),
	X845 => adc_samples(8459 DOWNTO 8450),
	X846 => adc_samples(8469 DOWNTO 8460),
	X847 => adc_samples(8479 DOWNTO 8470),
	X848 => adc_samples(8489 DOWNTO 8480),
	X849 => adc_samples(8499 DOWNTO 8490),
	X850 => adc_samples(8509 DOWNTO 8500),
	X851 => adc_samples(8519 DOWNTO 8510),
	X852 => adc_samples(8529 DOWNTO 8520),
	X853 => adc_samples(8539 DOWNTO 8530),
	X854 => adc_samples(8549 DOWNTO 8540),
	X855 => adc_samples(8559 DOWNTO 8550),
	X856 => adc_samples(8569 DOWNTO 8560),
	X857 => adc_samples(8579 DOWNTO 8570),
	X858 => adc_samples(8589 DOWNTO 8580),
	X859 => adc_samples(8599 DOWNTO 8590),
	X860 => adc_samples(8609 DOWNTO 8600),
	X861 => adc_samples(8619 DOWNTO 8610),
	X862 => adc_samples(8629 DOWNTO 8620),
	X863 => adc_samples(8639 DOWNTO 8630),
	X864 => adc_samples(8649 DOWNTO 8640),
	X865 => adc_samples(8659 DOWNTO 8650),
	X866 => adc_samples(8669 DOWNTO 8660),
	X867 => adc_samples(8679 DOWNTO 8670),
	X868 => adc_samples(8689 DOWNTO 8680),
	X869 => adc_samples(8699 DOWNTO 8690),
	X870 => adc_samples(8709 DOWNTO 8700),
	X871 => adc_samples(8719 DOWNTO 8710),
	X872 => adc_samples(8729 DOWNTO 8720),
	X873 => adc_samples(8739 DOWNTO 8730),
	X874 => adc_samples(8749 DOWNTO 8740),
	X875 => adc_samples(8759 DOWNTO 8750),
	X876 => adc_samples(8769 DOWNTO 8760),
	X877 => adc_samples(8779 DOWNTO 8770),
	X878 => adc_samples(8789 DOWNTO 8780),
	X879 => adc_samples(8799 DOWNTO 8790),
	X880 => adc_samples(8809 DOWNTO 8800),
	X881 => adc_samples(8819 DOWNTO 8810),
	X882 => adc_samples(8829 DOWNTO 8820),
	X883 => adc_samples(8839 DOWNTO 8830),
	X884 => adc_samples(8849 DOWNTO 8840),
	X885 => adc_samples(8859 DOWNTO 8850),
	X886 => adc_samples(8869 DOWNTO 8860),
	X887 => adc_samples(8879 DOWNTO 8870),
	X888 => adc_samples(8889 DOWNTO 8880),
	X889 => adc_samples(8899 DOWNTO 8890),
	X890 => adc_samples(8909 DOWNTO 8900),
	X891 => adc_samples(8919 DOWNTO 8910),
	X892 => adc_samples(8929 DOWNTO 8920),
	X893 => adc_samples(8939 DOWNTO 8930),
	X894 => adc_samples(8949 DOWNTO 8940),
	X895 => adc_samples(8959 DOWNTO 8950),
	X896 => adc_samples(8969 DOWNTO 8960),
	X897 => adc_samples(8979 DOWNTO 8970),
	X898 => adc_samples(8989 DOWNTO 8980),
	X899 => adc_samples(8999 DOWNTO 8990),
	X900 => adc_samples(9009 DOWNTO 9000),
	X901 => adc_samples(9019 DOWNTO 9010),
	X902 => adc_samples(9029 DOWNTO 9020),
	X903 => adc_samples(9039 DOWNTO 9030),
	X904 => adc_samples(9049 DOWNTO 9040),
	X905 => adc_samples(9059 DOWNTO 9050),
	X906 => adc_samples(9069 DOWNTO 9060),
	X907 => adc_samples(9079 DOWNTO 9070),
	X908 => adc_samples(9089 DOWNTO 9080),
	X909 => adc_samples(9099 DOWNTO 9090),
	X910 => adc_samples(9109 DOWNTO 9100),
	X911 => adc_samples(9119 DOWNTO 9110),
	X912 => adc_samples(9129 DOWNTO 9120),
	X913 => adc_samples(9139 DOWNTO 9130),
	X914 => adc_samples(9149 DOWNTO 9140),
	X915 => adc_samples(9159 DOWNTO 9150),
	X916 => adc_samples(9169 DOWNTO 9160),
	X917 => adc_samples(9179 DOWNTO 9170),
	X918 => adc_samples(9189 DOWNTO 9180),
	X919 => adc_samples(9199 DOWNTO 9190),
	X920 => adc_samples(9209 DOWNTO 9200),
	X921 => adc_samples(9219 DOWNTO 9210),
	X922 => adc_samples(9229 DOWNTO 9220),
	X923 => adc_samples(9239 DOWNTO 9230),
	X924 => adc_samples(9249 DOWNTO 9240),
	X925 => adc_samples(9259 DOWNTO 9250),
	X926 => adc_samples(9269 DOWNTO 9260),
	X927 => adc_samples(9279 DOWNTO 9270),
	X928 => adc_samples(9289 DOWNTO 9280),
	X929 => adc_samples(9299 DOWNTO 9290),
	X930 => adc_samples(9309 DOWNTO 9300),
	X931 => adc_samples(9319 DOWNTO 9310),
	X932 => adc_samples(9329 DOWNTO 9320),
	X933 => adc_samples(9339 DOWNTO 9330),
	X934 => adc_samples(9349 DOWNTO 9340),
	X935 => adc_samples(9359 DOWNTO 9350),
	X936 => adc_samples(9369 DOWNTO 9360),
	X937 => adc_samples(9379 DOWNTO 9370),
	X938 => adc_samples(9389 DOWNTO 9380),
	X939 => adc_samples(9399 DOWNTO 9390),
	X940 => adc_samples(9409 DOWNTO 9400),
	X941 => adc_samples(9419 DOWNTO 9410),
	X942 => adc_samples(9429 DOWNTO 9420),
	X943 => adc_samples(9439 DOWNTO 9430),
	X944 => adc_samples(9449 DOWNTO 9440),
	X945 => adc_samples(9459 DOWNTO 9450),
	X946 => adc_samples(9469 DOWNTO 9460),
	X947 => adc_samples(9479 DOWNTO 9470),
	X948 => adc_samples(9489 DOWNTO 9480),
	X949 => adc_samples(9499 DOWNTO 9490),
	X950 => adc_samples(9509 DOWNTO 9500),
	X951 => adc_samples(9519 DOWNTO 9510),
	X952 => adc_samples(9529 DOWNTO 9520),
	X953 => adc_samples(9539 DOWNTO 9530),
	X954 => adc_samples(9549 DOWNTO 9540),
	X955 => adc_samples(9559 DOWNTO 9550),
	X956 => adc_samples(9569 DOWNTO 9560),
	X957 => adc_samples(9579 DOWNTO 9570),
	X958 => adc_samples(9589 DOWNTO 9580),
	X959 => adc_samples(9599 DOWNTO 9590),
	X960 => adc_samples(9609 DOWNTO 9600),
	X961 => adc_samples(9619 DOWNTO 9610),
	X962 => adc_samples(9629 DOWNTO 9620),
	X963 => adc_samples(9639 DOWNTO 9630),
	X964 => adc_samples(9649 DOWNTO 9640),
	X965 => adc_samples(9659 DOWNTO 9650),
	X966 => adc_samples(9669 DOWNTO 9660),
	X967 => adc_samples(9679 DOWNTO 9670),
	X968 => adc_samples(9689 DOWNTO 9680),
	X969 => adc_samples(9699 DOWNTO 9690),
	X970 => adc_samples(9709 DOWNTO 9700),
	X971 => adc_samples(9719 DOWNTO 9710),
	X972 => adc_samples(9729 DOWNTO 9720),
	X973 => adc_samples(9739 DOWNTO 9730),
	X974 => adc_samples(9749 DOWNTO 9740),
	X975 => adc_samples(9759 DOWNTO 9750),
	X976 => adc_samples(9769 DOWNTO 9760),
	X977 => adc_samples(9779 DOWNTO 9770),
	X978 => adc_samples(9789 DOWNTO 9780),
	X979 => adc_samples(9799 DOWNTO 9790),
	X980 => adc_samples(9809 DOWNTO 9800),
	X981 => adc_samples(9819 DOWNTO 9810),
	X982 => adc_samples(9829 DOWNTO 9820),
	X983 => adc_samples(9839 DOWNTO 9830),
	X984 => adc_samples(9849 DOWNTO 9840),
	X985 => adc_samples(9859 DOWNTO 9850),
	X986 => adc_samples(9869 DOWNTO 9860),
	X987 => adc_samples(9879 DOWNTO 9870),
	X988 => adc_samples(9889 DOWNTO 9880),
	X989 => adc_samples(9899 DOWNTO 9890),
	X990 => adc_samples(9909 DOWNTO 9900),
	X991 => adc_samples(9919 DOWNTO 9910),
	X992 => adc_samples(9929 DOWNTO 9920),
	X993 => adc_samples(9939 DOWNTO 9930),
	X994 => adc_samples(9949 DOWNTO 9940),
	X995 => adc_samples(9959 DOWNTO 9950),
	X996 => adc_samples(9969 DOWNTO 9960),
	X997 => adc_samples(9979 DOWNTO 9970),
	X998 => adc_samples(9989 DOWNTO 9980),
	X999 => adc_samples(9999 DOWNTO 9990),
	X1000 => adc_samples(10009 DOWNTO 10000),
	X1001 => adc_samples(10019 DOWNTO 10010),
	X1002 => adc_samples(10029 DOWNTO 10020),
	X1003 => adc_samples(10039 DOWNTO 10030),
	X1004 => adc_samples(10049 DOWNTO 10040),
	X1005 => adc_samples(10059 DOWNTO 10050),
	X1006 => adc_samples(10069 DOWNTO 10060),
	X1007 => adc_samples(10079 DOWNTO 10070),
	X1008 => adc_samples(10089 DOWNTO 10080),
	X1009 => adc_samples(10099 DOWNTO 10090),
	X1010 => adc_samples(10109 DOWNTO 10100),
	X1011 => adc_samples(10119 DOWNTO 10110),
	X1012 => adc_samples(10129 DOWNTO 10120),
	X1013 => adc_samples(10139 DOWNTO 10130),
	X1014 => adc_samples(10149 DOWNTO 10140),
	X1015 => adc_samples(10159 DOWNTO 10150),
	X1016 => adc_samples(10169 DOWNTO 10160),
	X1017 => adc_samples(10179 DOWNTO 10170),
	X1018 => adc_samples(10189 DOWNTO 10180),
	X1019 => adc_samples(10199 DOWNTO 10190),
	X1020 => adc_samples(10209 DOWNTO 10200),
	X1021 => adc_samples(10219 DOWNTO 10210),
	X1022 => adc_samples(10229 DOWNTO 10220),
	X1023 => adc_samples(10239 DOWNTO 10230),
	X1024 => adc_samples(10249 DOWNTO 10240),
	X1025 => adc_samples(10259 DOWNTO 10250),
	X1026 => adc_samples(10269 DOWNTO 10260),
	X1027 => adc_samples(10279 DOWNTO 10270),
	X1028 => adc_samples(10289 DOWNTO 10280),
	X1029 => adc_samples(10299 DOWNTO 10290),
	X1030 => adc_samples(10309 DOWNTO 10300),
	X1031 => adc_samples(10319 DOWNTO 10310),
	X1032 => adc_samples(10329 DOWNTO 10320),
	X1033 => adc_samples(10339 DOWNTO 10330),
	X1034 => adc_samples(10349 DOWNTO 10340),
	X1035 => adc_samples(10359 DOWNTO 10350),
	X1036 => adc_samples(10369 DOWNTO 10360),
	X1037 => adc_samples(10379 DOWNTO 10370),
	X1038 => adc_samples(10389 DOWNTO 10380),
	X1039 => adc_samples(10399 DOWNTO 10390),
	X1040 => adc_samples(10409 DOWNTO 10400),
	X1041 => adc_samples(10419 DOWNTO 10410),
	X1042 => adc_samples(10429 DOWNTO 10420),
	X1043 => adc_samples(10439 DOWNTO 10430),
	X1044 => adc_samples(10449 DOWNTO 10440),
	X1045 => adc_samples(10459 DOWNTO 10450),
	X1046 => adc_samples(10469 DOWNTO 10460),
	X1047 => adc_samples(10479 DOWNTO 10470),
	X1048 => adc_samples(10489 DOWNTO 10480),
	X1049 => adc_samples(10499 DOWNTO 10490),
	X1050 => adc_samples(10509 DOWNTO 10500),
	X1051 => adc_samples(10519 DOWNTO 10510),
	X1052 => adc_samples(10529 DOWNTO 10520),
	X1053 => adc_samples(10539 DOWNTO 10530),
	X1054 => adc_samples(10549 DOWNTO 10540),
	X1055 => adc_samples(10559 DOWNTO 10550),
	X1056 => adc_samples(10569 DOWNTO 10560),
	X1057 => adc_samples(10579 DOWNTO 10570),
	X1058 => adc_samples(10589 DOWNTO 10580),
	X1059 => adc_samples(10599 DOWNTO 10590),
	X1060 => adc_samples(10609 DOWNTO 10600),
	X1061 => adc_samples(10619 DOWNTO 10610),
	X1062 => adc_samples(10629 DOWNTO 10620),
	X1063 => adc_samples(10639 DOWNTO 10630),
	X1064 => adc_samples(10649 DOWNTO 10640),
	X1065 => adc_samples(10659 DOWNTO 10650),
	X1066 => adc_samples(10669 DOWNTO 10660),
	X1067 => adc_samples(10679 DOWNTO 10670),
	X1068 => adc_samples(10689 DOWNTO 10680),
	X1069 => adc_samples(10699 DOWNTO 10690),
	X1070 => adc_samples(10709 DOWNTO 10700),
	X1071 => adc_samples(10719 DOWNTO 10710),
	X1072 => adc_samples(10729 DOWNTO 10720),
	X1073 => adc_samples(10739 DOWNTO 10730),
	X1074 => adc_samples(10749 DOWNTO 10740),
	X1075 => adc_samples(10759 DOWNTO 10750),
	X1076 => adc_samples(10769 DOWNTO 10760),
	X1077 => adc_samples(10779 DOWNTO 10770),
	X1078 => adc_samples(10789 DOWNTO 10780),
	X1079 => adc_samples(10799 DOWNTO 10790),
	X1080 => adc_samples(10809 DOWNTO 10800),
	X1081 => adc_samples(10819 DOWNTO 10810),
	X1082 => adc_samples(10829 DOWNTO 10820),
	X1083 => adc_samples(10839 DOWNTO 10830),
	X1084 => adc_samples(10849 DOWNTO 10840),
	X1085 => adc_samples(10859 DOWNTO 10850),
	X1086 => adc_samples(10869 DOWNTO 10860),
	X1087 => adc_samples(10879 DOWNTO 10870),
	X1088 => adc_samples(10889 DOWNTO 10880),
	X1089 => adc_samples(10899 DOWNTO 10890),
	X1090 => adc_samples(10909 DOWNTO 10900),
	X1091 => adc_samples(10919 DOWNTO 10910),
	X1092 => adc_samples(10929 DOWNTO 10920),
	X1093 => adc_samples(10939 DOWNTO 10930),
	X1094 => adc_samples(10949 DOWNTO 10940),
	X1095 => adc_samples(10959 DOWNTO 10950),
	X1096 => adc_samples(10969 DOWNTO 10960),
	X1097 => adc_samples(10979 DOWNTO 10970),
	X1098 => adc_samples(10989 DOWNTO 10980),
	X1099 => adc_samples(10999 DOWNTO 10990),
	X1100 => adc_samples(11009 DOWNTO 11000),
	X1101 => adc_samples(11019 DOWNTO 11010),
	X1102 => adc_samples(11029 DOWNTO 11020),
	X1103 => adc_samples(11039 DOWNTO 11030),
	X1104 => adc_samples(11049 DOWNTO 11040),
	X1105 => adc_samples(11059 DOWNTO 11050),
	X1106 => adc_samples(11069 DOWNTO 11060),
	X1107 => adc_samples(11079 DOWNTO 11070),
	X1108 => adc_samples(11089 DOWNTO 11080),
	X1109 => adc_samples(11099 DOWNTO 11090),
	X1110 => adc_samples(11109 DOWNTO 11100),
	X1111 => adc_samples(11119 DOWNTO 11110),
	X1112 => adc_samples(11129 DOWNTO 11120),
	X1113 => adc_samples(11139 DOWNTO 11130),
	X1114 => adc_samples(11149 DOWNTO 11140),
	X1115 => adc_samples(11159 DOWNTO 11150),
	X1116 => adc_samples(11169 DOWNTO 11160),
	X1117 => adc_samples(11179 DOWNTO 11170),
	X1118 => adc_samples(11189 DOWNTO 11180),
	X1119 => adc_samples(11199 DOWNTO 11190),
	X1120 => adc_samples(11209 DOWNTO 11200),
	X1121 => adc_samples(11219 DOWNTO 11210),
	X1122 => adc_samples(11229 DOWNTO 11220),
	X1123 => adc_samples(11239 DOWNTO 11230),
	X1124 => adc_samples(11249 DOWNTO 11240),
	X1125 => adc_samples(11259 DOWNTO 11250),
	X1126 => adc_samples(11269 DOWNTO 11260),
	X1127 => adc_samples(11279 DOWNTO 11270),
	X1128 => adc_samples(11289 DOWNTO 11280),
	X1129 => adc_samples(11299 DOWNTO 11290),
	X1130 => adc_samples(11309 DOWNTO 11300),
	X1131 => adc_samples(11319 DOWNTO 11310),
	X1132 => adc_samples(11329 DOWNTO 11320),
	X1133 => adc_samples(11339 DOWNTO 11330),
	X1134 => adc_samples(11349 DOWNTO 11340),
	X1135 => adc_samples(11359 DOWNTO 11350),
	X1136 => adc_samples(11369 DOWNTO 11360),
	X1137 => adc_samples(11379 DOWNTO 11370),
	X1138 => adc_samples(11389 DOWNTO 11380),
	X1139 => adc_samples(11399 DOWNTO 11390),
	X1140 => adc_samples(11409 DOWNTO 11400),
	X1141 => adc_samples(11419 DOWNTO 11410),
	X1142 => adc_samples(11429 DOWNTO 11420),
	X1143 => adc_samples(11439 DOWNTO 11430),
	X1144 => adc_samples(11449 DOWNTO 11440),
	X1145 => adc_samples(11459 DOWNTO 11450),
	X1146 => adc_samples(11469 DOWNTO 11460),
	X1147 => adc_samples(11479 DOWNTO 11470),
	X1148 => adc_samples(11489 DOWNTO 11480),
	X1149 => adc_samples(11499 DOWNTO 11490),
	X1150 => adc_samples(11509 DOWNTO 11500),
	X1151 => adc_samples(11519 DOWNTO 11510),
	X1152 => adc_samples(11529 DOWNTO 11520),
	X1153 => adc_samples(11539 DOWNTO 11530),
	X1154 => adc_samples(11549 DOWNTO 11540),
	X1155 => adc_samples(11559 DOWNTO 11550),
	X1156 => adc_samples(11569 DOWNTO 11560),
	X1157 => adc_samples(11579 DOWNTO 11570),
	X1158 => adc_samples(11589 DOWNTO 11580),
	X1159 => adc_samples(11599 DOWNTO 11590),
	X1160 => adc_samples(11609 DOWNTO 11600),
	X1161 => adc_samples(11619 DOWNTO 11610),
	X1162 => adc_samples(11629 DOWNTO 11620),
	X1163 => adc_samples(11639 DOWNTO 11630),
	X1164 => adc_samples(11649 DOWNTO 11640),
	X1165 => adc_samples(11659 DOWNTO 11650),
	X1166 => adc_samples(11669 DOWNTO 11660),
	X1167 => adc_samples(11679 DOWNTO 11670),
	X1168 => adc_samples(11689 DOWNTO 11680),
	X1169 => adc_samples(11699 DOWNTO 11690),
	X1170 => adc_samples(11709 DOWNTO 11700),
	X1171 => adc_samples(11719 DOWNTO 11710),
	X1172 => adc_samples(11729 DOWNTO 11720),
	X1173 => adc_samples(11739 DOWNTO 11730),
	X1174 => adc_samples(11749 DOWNTO 11740),
	X1175 => adc_samples(11759 DOWNTO 11750),
	X1176 => adc_samples(11769 DOWNTO 11760),
	X1177 => adc_samples(11779 DOWNTO 11770),
	X1178 => adc_samples(11789 DOWNTO 11780),
	X1179 => adc_samples(11799 DOWNTO 11790),
	X1180 => adc_samples(11809 DOWNTO 11800),
	X1181 => adc_samples(11819 DOWNTO 11810),
	X1182 => adc_samples(11829 DOWNTO 11820),
	X1183 => adc_samples(11839 DOWNTO 11830),
	X1184 => adc_samples(11849 DOWNTO 11840),
	X1185 => adc_samples(11859 DOWNTO 11850),
	X1186 => adc_samples(11869 DOWNTO 11860),
	X1187 => adc_samples(11879 DOWNTO 11870),
	X1188 => adc_samples(11889 DOWNTO 11880),
	X1189 => adc_samples(11899 DOWNTO 11890),
	X1190 => adc_samples(11909 DOWNTO 11900),
	X1191 => adc_samples(11919 DOWNTO 11910),
	X1192 => adc_samples(11929 DOWNTO 11920),
	X1193 => adc_samples(11939 DOWNTO 11930),
	X1194 => adc_samples(11949 DOWNTO 11940),
	X1195 => adc_samples(11959 DOWNTO 11950),
	X1196 => adc_samples(11969 DOWNTO 11960),
	X1197 => adc_samples(11979 DOWNTO 11970),
	X1198 => adc_samples(11989 DOWNTO 11980),
	X1199 => adc_samples(11999 DOWNTO 11990),
	X1200 => adc_samples(12009 DOWNTO 12000),
	X1201 => adc_samples(12019 DOWNTO 12010),
	X1202 => adc_samples(12029 DOWNTO 12020),
	X1203 => adc_samples(12039 DOWNTO 12030),
	X1204 => adc_samples(12049 DOWNTO 12040),
	X1205 => adc_samples(12059 DOWNTO 12050),
	X1206 => adc_samples(12069 DOWNTO 12060),
	X1207 => adc_samples(12079 DOWNTO 12070),
	X1208 => adc_samples(12089 DOWNTO 12080),
	X1209 => adc_samples(12099 DOWNTO 12090),
	X1210 => adc_samples(12109 DOWNTO 12100),
	X1211 => adc_samples(12119 DOWNTO 12110),
	X1212 => adc_samples(12129 DOWNTO 12120),
	X1213 => adc_samples(12139 DOWNTO 12130),
	X1214 => adc_samples(12149 DOWNTO 12140),
	X1215 => adc_samples(12159 DOWNTO 12150),
	X1216 => adc_samples(12169 DOWNTO 12160),
	X1217 => adc_samples(12179 DOWNTO 12170),
	X1218 => adc_samples(12189 DOWNTO 12180),
	X1219 => adc_samples(12199 DOWNTO 12190),
	X1220 => adc_samples(12209 DOWNTO 12200),
	X1221 => adc_samples(12219 DOWNTO 12210),
	X1222 => adc_samples(12229 DOWNTO 12220),
	X1223 => adc_samples(12239 DOWNTO 12230),
	X1224 => adc_samples(12249 DOWNTO 12240),
	X1225 => adc_samples(12259 DOWNTO 12250),
	X1226 => adc_samples(12269 DOWNTO 12260),
	X1227 => adc_samples(12279 DOWNTO 12270),
	X1228 => adc_samples(12289 DOWNTO 12280),
	X1229 => adc_samples(12299 DOWNTO 12290),
	X1230 => adc_samples(12309 DOWNTO 12300),
	X1231 => adc_samples(12319 DOWNTO 12310),
	X1232 => adc_samples(12329 DOWNTO 12320),
	X1233 => adc_samples(12339 DOWNTO 12330),
	X1234 => adc_samples(12349 DOWNTO 12340),
	X1235 => adc_samples(12359 DOWNTO 12350),
	X1236 => adc_samples(12369 DOWNTO 12360),
	X1237 => adc_samples(12379 DOWNTO 12370),
	X1238 => adc_samples(12389 DOWNTO 12380),
	X1239 => adc_samples(12399 DOWNTO 12390),
	X1240 => adc_samples(12409 DOWNTO 12400),
	X1241 => adc_samples(12419 DOWNTO 12410),
	X1242 => adc_samples(12429 DOWNTO 12420),
	X1243 => adc_samples(12439 DOWNTO 12430),
	X1244 => adc_samples(12449 DOWNTO 12440),
	X1245 => adc_samples(12459 DOWNTO 12450),
	X1246 => adc_samples(12469 DOWNTO 12460),
	X1247 => adc_samples(12479 DOWNTO 12470),
	X1248 => adc_samples(12489 DOWNTO 12480),
	X1249 => adc_samples(12499 DOWNTO 12490),
	X1250 => adc_samples(12509 DOWNTO 12500),
	X1251 => adc_samples(12519 DOWNTO 12510),
	X1252 => adc_samples(12529 DOWNTO 12520),
	X1253 => adc_samples(12539 DOWNTO 12530),
	X1254 => adc_samples(12549 DOWNTO 12540),
	X1255 => adc_samples(12559 DOWNTO 12550),
	X1256 => adc_samples(12569 DOWNTO 12560),
	X1257 => adc_samples(12579 DOWNTO 12570),
	X1258 => adc_samples(12589 DOWNTO 12580),
	X1259 => adc_samples(12599 DOWNTO 12590),
	X1260 => adc_samples(12609 DOWNTO 12600),
	X1261 => adc_samples(12619 DOWNTO 12610),
	X1262 => adc_samples(12629 DOWNTO 12620),
	X1263 => adc_samples(12639 DOWNTO 12630),
	X1264 => adc_samples(12649 DOWNTO 12640),
	X1265 => adc_samples(12659 DOWNTO 12650),
	X1266 => adc_samples(12669 DOWNTO 12660),
	X1267 => adc_samples(12679 DOWNTO 12670),
	X1268 => adc_samples(12689 DOWNTO 12680),
	X1269 => adc_samples(12699 DOWNTO 12690),
	X1270 => adc_samples(12709 DOWNTO 12700),
	X1271 => adc_samples(12719 DOWNTO 12710),
	X1272 => adc_samples(12729 DOWNTO 12720),
	X1273 => adc_samples(12739 DOWNTO 12730),
	X1274 => adc_samples(12749 DOWNTO 12740),
	X1275 => adc_samples(12759 DOWNTO 12750),
	X1276 => adc_samples(12769 DOWNTO 12760),
	X1277 => adc_samples(12779 DOWNTO 12770),
	X1278 => adc_samples(12789 DOWNTO 12780),
	X1279 => adc_samples(12799 DOWNTO 12790),
	X1280 => adc_samples(12809 DOWNTO 12800),
	X1281 => adc_samples(12819 DOWNTO 12810),
	X1282 => adc_samples(12829 DOWNTO 12820),
	X1283 => adc_samples(12839 DOWNTO 12830),
	X1284 => adc_samples(12849 DOWNTO 12840),
	X1285 => adc_samples(12859 DOWNTO 12850),
	X1286 => adc_samples(12869 DOWNTO 12860),
	X1287 => adc_samples(12879 DOWNTO 12870),
	X1288 => adc_samples(12889 DOWNTO 12880),
	X1289 => adc_samples(12899 DOWNTO 12890),
	X1290 => adc_samples(12909 DOWNTO 12900),
	X1291 => adc_samples(12919 DOWNTO 12910),
	X1292 => adc_samples(12929 DOWNTO 12920),
	X1293 => adc_samples(12939 DOWNTO 12930),
	X1294 => adc_samples(12949 DOWNTO 12940),
	X1295 => adc_samples(12959 DOWNTO 12950),
	X1296 => adc_samples(12969 DOWNTO 12960),
	X1297 => adc_samples(12979 DOWNTO 12970),
	X1298 => adc_samples(12989 DOWNTO 12980),
	X1299 => adc_samples(12999 DOWNTO 12990),
	X1300 => adc_samples(13009 DOWNTO 13000),
	X1301 => adc_samples(13019 DOWNTO 13010),
	X1302 => adc_samples(13029 DOWNTO 13020),
	X1303 => adc_samples(13039 DOWNTO 13030),
	X1304 => adc_samples(13049 DOWNTO 13040),
	X1305 => adc_samples(13059 DOWNTO 13050),
	X1306 => adc_samples(13069 DOWNTO 13060),
	X1307 => adc_samples(13079 DOWNTO 13070),
	X1308 => adc_samples(13089 DOWNTO 13080),
	X1309 => adc_samples(13099 DOWNTO 13090),
	X1310 => adc_samples(13109 DOWNTO 13100),
	X1311 => adc_samples(13119 DOWNTO 13110),
	X1312 => adc_samples(13129 DOWNTO 13120),
	X1313 => adc_samples(13139 DOWNTO 13130),
	X1314 => adc_samples(13149 DOWNTO 13140),
	X1315 => adc_samples(13159 DOWNTO 13150),
	X1316 => adc_samples(13169 DOWNTO 13160),
	X1317 => adc_samples(13179 DOWNTO 13170),
	X1318 => adc_samples(13189 DOWNTO 13180),
	X1319 => adc_samples(13199 DOWNTO 13190),
	X1320 => adc_samples(13209 DOWNTO 13200),
	X1321 => adc_samples(13219 DOWNTO 13210),
	X1322 => adc_samples(13229 DOWNTO 13220),
	X1323 => adc_samples(13239 DOWNTO 13230),
	X1324 => adc_samples(13249 DOWNTO 13240),
	X1325 => adc_samples(13259 DOWNTO 13250),
	X1326 => adc_samples(13269 DOWNTO 13260),
	X1327 => adc_samples(13279 DOWNTO 13270),
	X1328 => adc_samples(13289 DOWNTO 13280),
	X1329 => adc_samples(13299 DOWNTO 13290),
	X1330 => adc_samples(13309 DOWNTO 13300),
	X1331 => adc_samples(13319 DOWNTO 13310),
	X1332 => adc_samples(13329 DOWNTO 13320),
	X1333 => adc_samples(13339 DOWNTO 13330),
	X1334 => adc_samples(13349 DOWNTO 13340),
	X1335 => adc_samples(13359 DOWNTO 13350),
	X1336 => adc_samples(13369 DOWNTO 13360),
	X1337 => adc_samples(13379 DOWNTO 13370),
	X1338 => adc_samples(13389 DOWNTO 13380),
	X1339 => adc_samples(13399 DOWNTO 13390),
	X1340 => adc_samples(13409 DOWNTO 13400),
	X1341 => adc_samples(13419 DOWNTO 13410),
	X1342 => adc_samples(13429 DOWNTO 13420),
	X1343 => adc_samples(13439 DOWNTO 13430),
	X1344 => adc_samples(13449 DOWNTO 13440),
	X1345 => adc_samples(13459 DOWNTO 13450),
	X1346 => adc_samples(13469 DOWNTO 13460),
	X1347 => adc_samples(13479 DOWNTO 13470),
	X1348 => adc_samples(13489 DOWNTO 13480),
	X1349 => adc_samples(13499 DOWNTO 13490),
	X1350 => adc_samples(13509 DOWNTO 13500),
	X1351 => adc_samples(13519 DOWNTO 13510),
	X1352 => adc_samples(13529 DOWNTO 13520),
	X1353 => adc_samples(13539 DOWNTO 13530),
	X1354 => adc_samples(13549 DOWNTO 13540),
	X1355 => adc_samples(13559 DOWNTO 13550),
	X1356 => adc_samples(13569 DOWNTO 13560),
	X1357 => adc_samples(13579 DOWNTO 13570),
	X1358 => adc_samples(13589 DOWNTO 13580),
	X1359 => adc_samples(13599 DOWNTO 13590),
	X1360 => adc_samples(13609 DOWNTO 13600),
	X1361 => adc_samples(13619 DOWNTO 13610),
	X1362 => adc_samples(13629 DOWNTO 13620),
	X1363 => adc_samples(13639 DOWNTO 13630),
	X1364 => adc_samples(13649 DOWNTO 13640),
	X1365 => adc_samples(13659 DOWNTO 13650),
	X1366 => adc_samples(13669 DOWNTO 13660),
	X1367 => adc_samples(13679 DOWNTO 13670),
	X1368 => adc_samples(13689 DOWNTO 13680),
	X1369 => adc_samples(13699 DOWNTO 13690),
	X1370 => adc_samples(13709 DOWNTO 13700),
	X1371 => adc_samples(13719 DOWNTO 13710),
	X1372 => adc_samples(13729 DOWNTO 13720),
	X1373 => adc_samples(13739 DOWNTO 13730),
	X1374 => adc_samples(13749 DOWNTO 13740),
	X1375 => adc_samples(13759 DOWNTO 13750),
	X1376 => adc_samples(13769 DOWNTO 13760),
	X1377 => adc_samples(13779 DOWNTO 13770),
	X1378 => adc_samples(13789 DOWNTO 13780),
	X1379 => adc_samples(13799 DOWNTO 13790),
	X1380 => adc_samples(13809 DOWNTO 13800),
	X1381 => adc_samples(13819 DOWNTO 13810),
	X1382 => adc_samples(13829 DOWNTO 13820),
	X1383 => adc_samples(13839 DOWNTO 13830),
	X1384 => adc_samples(13849 DOWNTO 13840),
	X1385 => adc_samples(13859 DOWNTO 13850),
	X1386 => adc_samples(13869 DOWNTO 13860),
	X1387 => adc_samples(13879 DOWNTO 13870),
	X1388 => adc_samples(13889 DOWNTO 13880),
	X1389 => adc_samples(13899 DOWNTO 13890),
	X1390 => adc_samples(13909 DOWNTO 13900),
	X1391 => adc_samples(13919 DOWNTO 13910),
	X1392 => adc_samples(13929 DOWNTO 13920),
	X1393 => adc_samples(13939 DOWNTO 13930),
	X1394 => adc_samples(13949 DOWNTO 13940),
	X1395 => adc_samples(13959 DOWNTO 13950),
	X1396 => adc_samples(13969 DOWNTO 13960),
	X1397 => adc_samples(13979 DOWNTO 13970),
	X1398 => adc_samples(13989 DOWNTO 13980),
	X1399 => adc_samples(13999 DOWNTO 13990),
	X1400 => adc_samples(14009 DOWNTO 14000),
	X1401 => adc_samples(14019 DOWNTO 14010),
	X1402 => adc_samples(14029 DOWNTO 14020),
	X1403 => adc_samples(14039 DOWNTO 14030),
	X1404 => adc_samples(14049 DOWNTO 14040),
	X1405 => adc_samples(14059 DOWNTO 14050),
	X1406 => adc_samples(14069 DOWNTO 14060),
	X1407 => adc_samples(14079 DOWNTO 14070),
	X1408 => adc_samples(14089 DOWNTO 14080),
	X1409 => adc_samples(14099 DOWNTO 14090),
	X1410 => adc_samples(14109 DOWNTO 14100),
	X1411 => adc_samples(14119 DOWNTO 14110),
	X1412 => adc_samples(14129 DOWNTO 14120),
	X1413 => adc_samples(14139 DOWNTO 14130),
	X1414 => adc_samples(14149 DOWNTO 14140),
	X1415 => adc_samples(14159 DOWNTO 14150),
	X1416 => adc_samples(14169 DOWNTO 14160),
	X1417 => adc_samples(14179 DOWNTO 14170),
	X1418 => adc_samples(14189 DOWNTO 14180),
	X1419 => adc_samples(14199 DOWNTO 14190),
	X1420 => adc_samples(14209 DOWNTO 14200),
	X1421 => adc_samples(14219 DOWNTO 14210),
	X1422 => adc_samples(14229 DOWNTO 14220),
	X1423 => adc_samples(14239 DOWNTO 14230),
	X1424 => adc_samples(14249 DOWNTO 14240),
	X1425 => adc_samples(14259 DOWNTO 14250),
	X1426 => adc_samples(14269 DOWNTO 14260),
	X1427 => adc_samples(14279 DOWNTO 14270),
	X1428 => adc_samples(14289 DOWNTO 14280),
	X1429 => adc_samples(14299 DOWNTO 14290),
	X1430 => adc_samples(14309 DOWNTO 14300),
	X1431 => adc_samples(14319 DOWNTO 14310),
	X1432 => adc_samples(14329 DOWNTO 14320),
	X1433 => adc_samples(14339 DOWNTO 14330),
	X1434 => adc_samples(14349 DOWNTO 14340),
	X1435 => adc_samples(14359 DOWNTO 14350),
	X1436 => adc_samples(14369 DOWNTO 14360),
	X1437 => adc_samples(14379 DOWNTO 14370),
	X1438 => adc_samples(14389 DOWNTO 14380),
	X1439 => adc_samples(14399 DOWNTO 14390),
	X1440 => adc_samples(14409 DOWNTO 14400),
	X1441 => adc_samples(14419 DOWNTO 14410),
	X1442 => adc_samples(14429 DOWNTO 14420),
	X1443 => adc_samples(14439 DOWNTO 14430),
	X1444 => adc_samples(14449 DOWNTO 14440),
	X1445 => adc_samples(14459 DOWNTO 14450),
	X1446 => adc_samples(14469 DOWNTO 14460),
	X1447 => adc_samples(14479 DOWNTO 14470),
	X1448 => adc_samples(14489 DOWNTO 14480),
	X1449 => adc_samples(14499 DOWNTO 14490),
	X1450 => adc_samples(14509 DOWNTO 14500),
	X1451 => adc_samples(14519 DOWNTO 14510),
	X1452 => adc_samples(14529 DOWNTO 14520),
	X1453 => adc_samples(14539 DOWNTO 14530),
	X1454 => adc_samples(14549 DOWNTO 14540),
	X1455 => adc_samples(14559 DOWNTO 14550),
	X1456 => adc_samples(14569 DOWNTO 14560),
	X1457 => adc_samples(14579 DOWNTO 14570),
	X1458 => adc_samples(14589 DOWNTO 14580),
	X1459 => adc_samples(14599 DOWNTO 14590),
	X1460 => adc_samples(14609 DOWNTO 14600),
	X1461 => adc_samples(14619 DOWNTO 14610),
	X1462 => adc_samples(14629 DOWNTO 14620),
	X1463 => adc_samples(14639 DOWNTO 14630),
	X1464 => adc_samples(14649 DOWNTO 14640),
	X1465 => adc_samples(14659 DOWNTO 14650),
	X1466 => adc_samples(14669 DOWNTO 14660),
	X1467 => adc_samples(14679 DOWNTO 14670),
	X1468 => adc_samples(14689 DOWNTO 14680),
	X1469 => adc_samples(14699 DOWNTO 14690),
	X1470 => adc_samples(14709 DOWNTO 14700),
	X1471 => adc_samples(14719 DOWNTO 14710),
	X1472 => adc_samples(14729 DOWNTO 14720),
	X1473 => adc_samples(14739 DOWNTO 14730),
	X1474 => adc_samples(14749 DOWNTO 14740),
	X1475 => adc_samples(14759 DOWNTO 14750),
	X1476 => adc_samples(14769 DOWNTO 14760),
	X1477 => adc_samples(14779 DOWNTO 14770),
	X1478 => adc_samples(14789 DOWNTO 14780),
	X1479 => adc_samples(14799 DOWNTO 14790),
	X1480 => adc_samples(14809 DOWNTO 14800),
	X1481 => adc_samples(14819 DOWNTO 14810),
	X1482 => adc_samples(14829 DOWNTO 14820),
	X1483 => adc_samples(14839 DOWNTO 14830),
	X1484 => adc_samples(14849 DOWNTO 14840),
	X1485 => adc_samples(14859 DOWNTO 14850),
	X1486 => adc_samples(14869 DOWNTO 14860),
	X1487 => adc_samples(14879 DOWNTO 14870),
	X1488 => adc_samples(14889 DOWNTO 14880),
	X1489 => adc_samples(14899 DOWNTO 14890),
	X1490 => adc_samples(14909 DOWNTO 14900),
	X1491 => adc_samples(14919 DOWNTO 14910),
	X1492 => adc_samples(14929 DOWNTO 14920),
	X1493 => adc_samples(14939 DOWNTO 14930),
	X1494 => adc_samples(14949 DOWNTO 14940),
	X1495 => adc_samples(14959 DOWNTO 14950),
	X1496 => adc_samples(14969 DOWNTO 14960),
	X1497 => adc_samples(14979 DOWNTO 14970),
	X1498 => adc_samples(14989 DOWNTO 14980),
	X1499 => adc_samples(14999 DOWNTO 14990),
	X1500 => adc_samples(15009 DOWNTO 15000),
	X1501 => adc_samples(15019 DOWNTO 15010),
	X1502 => adc_samples(15029 DOWNTO 15020),
	X1503 => adc_samples(15039 DOWNTO 15030),
	X1504 => adc_samples(15049 DOWNTO 15040),
	X1505 => adc_samples(15059 DOWNTO 15050),
	X1506 => adc_samples(15069 DOWNTO 15060),
	X1507 => adc_samples(15079 DOWNTO 15070),
	X1508 => adc_samples(15089 DOWNTO 15080),
	X1509 => adc_samples(15099 DOWNTO 15090),
	X1510 => adc_samples(15109 DOWNTO 15100),
	X1511 => adc_samples(15119 DOWNTO 15110),
	X1512 => adc_samples(15129 DOWNTO 15120),
	X1513 => adc_samples(15139 DOWNTO 15130),
	X1514 => adc_samples(15149 DOWNTO 15140),
	X1515 => adc_samples(15159 DOWNTO 15150),
	X1516 => adc_samples(15169 DOWNTO 15160),
	X1517 => adc_samples(15179 DOWNTO 15170),
	X1518 => adc_samples(15189 DOWNTO 15180),
	X1519 => adc_samples(15199 DOWNTO 15190),
	X1520 => adc_samples(15209 DOWNTO 15200),
	X1521 => adc_samples(15219 DOWNTO 15210),
	X1522 => adc_samples(15229 DOWNTO 15220),
	X1523 => adc_samples(15239 DOWNTO 15230),
	X1524 => adc_samples(15249 DOWNTO 15240),
	X1525 => adc_samples(15259 DOWNTO 15250),
	X1526 => adc_samples(15269 DOWNTO 15260),
	X1527 => adc_samples(15279 DOWNTO 15270),
	X1528 => adc_samples(15289 DOWNTO 15280),
	X1529 => adc_samples(15299 DOWNTO 15290),
	X1530 => adc_samples(15309 DOWNTO 15300),
	X1531 => adc_samples(15319 DOWNTO 15310),
	X1532 => adc_samples(15329 DOWNTO 15320),
	X1533 => adc_samples(15339 DOWNTO 15330),
	X1534 => adc_samples(15349 DOWNTO 15340),
	X1535 => adc_samples(15359 DOWNTO 15350),
	X1536 => adc_samples(15369 DOWNTO 15360),
	X1537 => adc_samples(15379 DOWNTO 15370),
	X1538 => adc_samples(15389 DOWNTO 15380),
	X1539 => adc_samples(15399 DOWNTO 15390),
	X1540 => adc_samples(15409 DOWNTO 15400),
	X1541 => adc_samples(15419 DOWNTO 15410),
	X1542 => adc_samples(15429 DOWNTO 15420),
	X1543 => adc_samples(15439 DOWNTO 15430),
	X1544 => adc_samples(15449 DOWNTO 15440),
	X1545 => adc_samples(15459 DOWNTO 15450),
	X1546 => adc_samples(15469 DOWNTO 15460),
	X1547 => adc_samples(15479 DOWNTO 15470),
	X1548 => adc_samples(15489 DOWNTO 15480),
	X1549 => adc_samples(15499 DOWNTO 15490),
	X1550 => adc_samples(15509 DOWNTO 15500),
	X1551 => adc_samples(15519 DOWNTO 15510),
	X1552 => adc_samples(15529 DOWNTO 15520),
	X1553 => adc_samples(15539 DOWNTO 15530),
	X1554 => adc_samples(15549 DOWNTO 15540),
	X1555 => adc_samples(15559 DOWNTO 15550),
	X1556 => adc_samples(15569 DOWNTO 15560),
	X1557 => adc_samples(15579 DOWNTO 15570),
	X1558 => adc_samples(15589 DOWNTO 15580),
	X1559 => adc_samples(15599 DOWNTO 15590),
	X1560 => adc_samples(15609 DOWNTO 15600),
	X1561 => adc_samples(15619 DOWNTO 15610),
	X1562 => adc_samples(15629 DOWNTO 15620),
	X1563 => adc_samples(15639 DOWNTO 15630),
	X1564 => adc_samples(15649 DOWNTO 15640),
	X1565 => adc_samples(15659 DOWNTO 15650),
	X1566 => adc_samples(15669 DOWNTO 15660),
	X1567 => adc_samples(15679 DOWNTO 15670),
	X1568 => adc_samples(15689 DOWNTO 15680),
	X1569 => adc_samples(15699 DOWNTO 15690),
	X1570 => adc_samples(15709 DOWNTO 15700),
	X1571 => adc_samples(15719 DOWNTO 15710),
	X1572 => adc_samples(15729 DOWNTO 15720),
	X1573 => adc_samples(15739 DOWNTO 15730),
	X1574 => adc_samples(15749 DOWNTO 15740),
	X1575 => adc_samples(15759 DOWNTO 15750),
	X1576 => adc_samples(15769 DOWNTO 15760),
	X1577 => adc_samples(15779 DOWNTO 15770),
	X1578 => adc_samples(15789 DOWNTO 15780),
	X1579 => adc_samples(15799 DOWNTO 15790),
	X1580 => adc_samples(15809 DOWNTO 15800),
	X1581 => adc_samples(15819 DOWNTO 15810),
	X1582 => adc_samples(15829 DOWNTO 15820),
	X1583 => adc_samples(15839 DOWNTO 15830),
	X1584 => adc_samples(15849 DOWNTO 15840),
	X1585 => adc_samples(15859 DOWNTO 15850),
	X1586 => adc_samples(15869 DOWNTO 15860),
	X1587 => adc_samples(15879 DOWNTO 15870),
	X1588 => adc_samples(15889 DOWNTO 15880),
	X1589 => adc_samples(15899 DOWNTO 15890),
	X1590 => adc_samples(15909 DOWNTO 15900),
	X1591 => adc_samples(15919 DOWNTO 15910),
	X1592 => adc_samples(15929 DOWNTO 15920),
	X1593 => adc_samples(15939 DOWNTO 15930),
	X1594 => adc_samples(15949 DOWNTO 15940),
	X1595 => adc_samples(15959 DOWNTO 15950),
	X1596 => adc_samples(15969 DOWNTO 15960),
	X1597 => adc_samples(15979 DOWNTO 15970),
	X1598 => adc_samples(15989 DOWNTO 15980),
	X1599 => adc_samples(15999 DOWNTO 15990),
	X1600 => adc_samples(16009 DOWNTO 16000),
	X1601 => adc_samples(16019 DOWNTO 16010),
	X1602 => adc_samples(16029 DOWNTO 16020),
	X1603 => adc_samples(16039 DOWNTO 16030),
	X1604 => adc_samples(16049 DOWNTO 16040),
	X1605 => adc_samples(16059 DOWNTO 16050),
	X1606 => adc_samples(16069 DOWNTO 16060),
	X1607 => adc_samples(16079 DOWNTO 16070),
	X1608 => adc_samples(16089 DOWNTO 16080),
	X1609 => adc_samples(16099 DOWNTO 16090),
	X1610 => adc_samples(16109 DOWNTO 16100),
	X1611 => adc_samples(16119 DOWNTO 16110),
	X1612 => adc_samples(16129 DOWNTO 16120),
	X1613 => adc_samples(16139 DOWNTO 16130),
	X1614 => adc_samples(16149 DOWNTO 16140),
	X1615 => adc_samples(16159 DOWNTO 16150),
	X1616 => adc_samples(16169 DOWNTO 16160),
	X1617 => adc_samples(16179 DOWNTO 16170),
	X1618 => adc_samples(16189 DOWNTO 16180),
	X1619 => adc_samples(16199 DOWNTO 16190),
	X1620 => adc_samples(16209 DOWNTO 16200),
	X1621 => adc_samples(16219 DOWNTO 16210),
	X1622 => adc_samples(16229 DOWNTO 16220),
	X1623 => adc_samples(16239 DOWNTO 16230),
	X1624 => adc_samples(16249 DOWNTO 16240),
	X1625 => adc_samples(16259 DOWNTO 16250),
	X1626 => adc_samples(16269 DOWNTO 16260),
	X1627 => adc_samples(16279 DOWNTO 16270),
	X1628 => adc_samples(16289 DOWNTO 16280),
	X1629 => adc_samples(16299 DOWNTO 16290),
	X1630 => adc_samples(16309 DOWNTO 16300),
	X1631 => adc_samples(16319 DOWNTO 16310),
	X1632 => adc_samples(16329 DOWNTO 16320),
	X1633 => adc_samples(16339 DOWNTO 16330),
	X1634 => adc_samples(16349 DOWNTO 16340),
	X1635 => adc_samples(16359 DOWNTO 16350),
	X1636 => adc_samples(16369 DOWNTO 16360),
	X1637 => adc_samples(16379 DOWNTO 16370),
	X1638 => adc_samples(16389 DOWNTO 16380),
	X1639 => adc_samples(16399 DOWNTO 16390),
	X1640 => adc_samples(16409 DOWNTO 16400),
	X1641 => adc_samples(16419 DOWNTO 16410),
	X1642 => adc_samples(16429 DOWNTO 16420),
	X1643 => adc_samples(16439 DOWNTO 16430),
	X1644 => adc_samples(16449 DOWNTO 16440),
	X1645 => adc_samples(16459 DOWNTO 16450),
	X1646 => adc_samples(16469 DOWNTO 16460),
	X1647 => adc_samples(16479 DOWNTO 16470),
	X1648 => adc_samples(16489 DOWNTO 16480),
	X1649 => adc_samples(16499 DOWNTO 16490),
	X1650 => adc_samples(16509 DOWNTO 16500),
	X1651 => adc_samples(16519 DOWNTO 16510),
	X1652 => adc_samples(16529 DOWNTO 16520),
	X1653 => adc_samples(16539 DOWNTO 16530),
	X1654 => adc_samples(16549 DOWNTO 16540),
	X1655 => adc_samples(16559 DOWNTO 16550),
	X1656 => adc_samples(16569 DOWNTO 16560),
	X1657 => adc_samples(16579 DOWNTO 16570),
	X1658 => adc_samples(16589 DOWNTO 16580),
	X1659 => adc_samples(16599 DOWNTO 16590),
	X1660 => adc_samples(16609 DOWNTO 16600),
	X1661 => adc_samples(16619 DOWNTO 16610),
	X1662 => adc_samples(16629 DOWNTO 16620),
	X1663 => adc_samples(16639 DOWNTO 16630),
	X1664 => adc_samples(16649 DOWNTO 16640),
	X1665 => adc_samples(16659 DOWNTO 16650),
	X1666 => adc_samples(16669 DOWNTO 16660),
	X1667 => adc_samples(16679 DOWNTO 16670),
	X1668 => adc_samples(16689 DOWNTO 16680),
	X1669 => adc_samples(16699 DOWNTO 16690),
	X1670 => adc_samples(16709 DOWNTO 16700),
	X1671 => adc_samples(16719 DOWNTO 16710),
	X1672 => adc_samples(16729 DOWNTO 16720),
	X1673 => adc_samples(16739 DOWNTO 16730),
	X1674 => adc_samples(16749 DOWNTO 16740),
	X1675 => adc_samples(16759 DOWNTO 16750),
	X1676 => adc_samples(16769 DOWNTO 16760),
	X1677 => adc_samples(16779 DOWNTO 16770),
	X1678 => adc_samples(16789 DOWNTO 16780),
	X1679 => adc_samples(16799 DOWNTO 16790),
	X1680 => adc_samples(16809 DOWNTO 16800),
	X1681 => adc_samples(16819 DOWNTO 16810),
	X1682 => adc_samples(16829 DOWNTO 16820),
	X1683 => adc_samples(16839 DOWNTO 16830),
	X1684 => adc_samples(16849 DOWNTO 16840),
	X1685 => adc_samples(16859 DOWNTO 16850),
	X1686 => adc_samples(16869 DOWNTO 16860),
	X1687 => adc_samples(16879 DOWNTO 16870),
	X1688 => adc_samples(16889 DOWNTO 16880),
	X1689 => adc_samples(16899 DOWNTO 16890),
	X1690 => adc_samples(16909 DOWNTO 16900),
	X1691 => adc_samples(16919 DOWNTO 16910),
	X1692 => adc_samples(16929 DOWNTO 16920),
	X1693 => adc_samples(16939 DOWNTO 16930),
	X1694 => adc_samples(16949 DOWNTO 16940),
	X1695 => adc_samples(16959 DOWNTO 16950),
	X1696 => adc_samples(16969 DOWNTO 16960),
	X1697 => adc_samples(16979 DOWNTO 16970),
	X1698 => adc_samples(16989 DOWNTO 16980),
	X1699 => adc_samples(16999 DOWNTO 16990),
	X1700 => adc_samples(17009 DOWNTO 17000),
	X1701 => adc_samples(17019 DOWNTO 17010),
	X1702 => adc_samples(17029 DOWNTO 17020),
	X1703 => adc_samples(17039 DOWNTO 17030),
	X1704 => adc_samples(17049 DOWNTO 17040),
	X1705 => adc_samples(17059 DOWNTO 17050),
	X1706 => adc_samples(17069 DOWNTO 17060),
	X1707 => adc_samples(17079 DOWNTO 17070),
	X1708 => adc_samples(17089 DOWNTO 17080),
	X1709 => adc_samples(17099 DOWNTO 17090),
	X1710 => adc_samples(17109 DOWNTO 17100),
	X1711 => adc_samples(17119 DOWNTO 17110),
	X1712 => adc_samples(17129 DOWNTO 17120),
	X1713 => adc_samples(17139 DOWNTO 17130),
	X1714 => adc_samples(17149 DOWNTO 17140),
	X1715 => adc_samples(17159 DOWNTO 17150),
	X1716 => adc_samples(17169 DOWNTO 17160),
	X1717 => adc_samples(17179 DOWNTO 17170),
	X1718 => adc_samples(17189 DOWNTO 17180),
	X1719 => adc_samples(17199 DOWNTO 17190),
	X1720 => adc_samples(17209 DOWNTO 17200),
	X1721 => adc_samples(17219 DOWNTO 17210),
	X1722 => adc_samples(17229 DOWNTO 17220),
	X1723 => adc_samples(17239 DOWNTO 17230),
	X1724 => adc_samples(17249 DOWNTO 17240),
	X1725 => adc_samples(17259 DOWNTO 17250),
	X1726 => adc_samples(17269 DOWNTO 17260),
	X1727 => adc_samples(17279 DOWNTO 17270),
	X1728 => adc_samples(17289 DOWNTO 17280),
	X1729 => adc_samples(17299 DOWNTO 17290),
	X1730 => adc_samples(17309 DOWNTO 17300),
	X1731 => adc_samples(17319 DOWNTO 17310),
	X1732 => adc_samples(17329 DOWNTO 17320),
	X1733 => adc_samples(17339 DOWNTO 17330),
	X1734 => adc_samples(17349 DOWNTO 17340),
	X1735 => adc_samples(17359 DOWNTO 17350),
	X1736 => adc_samples(17369 DOWNTO 17360),
	X1737 => adc_samples(17379 DOWNTO 17370),
	X1738 => adc_samples(17389 DOWNTO 17380),
	X1739 => adc_samples(17399 DOWNTO 17390),
	X1740 => adc_samples(17409 DOWNTO 17400),
	X1741 => adc_samples(17419 DOWNTO 17410),
	X1742 => adc_samples(17429 DOWNTO 17420),
	X1743 => adc_samples(17439 DOWNTO 17430),
	X1744 => adc_samples(17449 DOWNTO 17440),
	X1745 => adc_samples(17459 DOWNTO 17450),
	X1746 => adc_samples(17469 DOWNTO 17460),
	X1747 => adc_samples(17479 DOWNTO 17470),
	X1748 => adc_samples(17489 DOWNTO 17480),
	X1749 => adc_samples(17499 DOWNTO 17490),
	X1750 => adc_samples(17509 DOWNTO 17500),
	X1751 => adc_samples(17519 DOWNTO 17510),
	X1752 => adc_samples(17529 DOWNTO 17520),
	X1753 => adc_samples(17539 DOWNTO 17530),
	X1754 => adc_samples(17549 DOWNTO 17540),
	X1755 => adc_samples(17559 DOWNTO 17550),
	X1756 => adc_samples(17569 DOWNTO 17560),
	X1757 => adc_samples(17579 DOWNTO 17570),
	X1758 => adc_samples(17589 DOWNTO 17580),
	X1759 => adc_samples(17599 DOWNTO 17590),
	X1760 => adc_samples(17609 DOWNTO 17600),
	X1761 => adc_samples(17619 DOWNTO 17610),
	X1762 => adc_samples(17629 DOWNTO 17620),
	X1763 => adc_samples(17639 DOWNTO 17630),
	X1764 => adc_samples(17649 DOWNTO 17640),
	X1765 => adc_samples(17659 DOWNTO 17650),
	X1766 => adc_samples(17669 DOWNTO 17660),
	X1767 => adc_samples(17679 DOWNTO 17670),
	X1768 => adc_samples(17689 DOWNTO 17680),
	X1769 => adc_samples(17699 DOWNTO 17690),
	X1770 => adc_samples(17709 DOWNTO 17700),
	X1771 => adc_samples(17719 DOWNTO 17710),
	X1772 => adc_samples(17729 DOWNTO 17720),
	X1773 => adc_samples(17739 DOWNTO 17730),
	X1774 => adc_samples(17749 DOWNTO 17740),
	X1775 => adc_samples(17759 DOWNTO 17750),
	X1776 => adc_samples(17769 DOWNTO 17760),
	X1777 => adc_samples(17779 DOWNTO 17770),
	X1778 => adc_samples(17789 DOWNTO 17780),
	X1779 => adc_samples(17799 DOWNTO 17790),
	X1780 => adc_samples(17809 DOWNTO 17800),
	X1781 => adc_samples(17819 DOWNTO 17810),
	X1782 => adc_samples(17829 DOWNTO 17820),
	X1783 => adc_samples(17839 DOWNTO 17830),
	X1784 => adc_samples(17849 DOWNTO 17840),
	X1785 => adc_samples(17859 DOWNTO 17850),
	X1786 => adc_samples(17869 DOWNTO 17860),
	X1787 => adc_samples(17879 DOWNTO 17870),
	X1788 => adc_samples(17889 DOWNTO 17880),
	X1789 => adc_samples(17899 DOWNTO 17890),
	X1790 => adc_samples(17909 DOWNTO 17900),
	X1791 => adc_samples(17919 DOWNTO 17910),
	X1792 => adc_samples(17929 DOWNTO 17920),
	X1793 => adc_samples(17939 DOWNTO 17930),
	X1794 => adc_samples(17949 DOWNTO 17940),
	X1795 => adc_samples(17959 DOWNTO 17950),
	X1796 => adc_samples(17969 DOWNTO 17960),
	X1797 => adc_samples(17979 DOWNTO 17970),
	X1798 => adc_samples(17989 DOWNTO 17980),
	X1799 => adc_samples(17999 DOWNTO 17990),
	X1800 => adc_samples(18009 DOWNTO 18000),
	X1801 => adc_samples(18019 DOWNTO 18010),
	X1802 => adc_samples(18029 DOWNTO 18020),
	X1803 => adc_samples(18039 DOWNTO 18030),
	X1804 => adc_samples(18049 DOWNTO 18040),
	X1805 => adc_samples(18059 DOWNTO 18050),
	X1806 => adc_samples(18069 DOWNTO 18060),
	X1807 => adc_samples(18079 DOWNTO 18070),
	X1808 => adc_samples(18089 DOWNTO 18080),
	X1809 => adc_samples(18099 DOWNTO 18090),
	X1810 => adc_samples(18109 DOWNTO 18100),
	X1811 => adc_samples(18119 DOWNTO 18110),
	X1812 => adc_samples(18129 DOWNTO 18120),
	X1813 => adc_samples(18139 DOWNTO 18130),
	X1814 => adc_samples(18149 DOWNTO 18140),
	X1815 => adc_samples(18159 DOWNTO 18150),
	X1816 => adc_samples(18169 DOWNTO 18160),
	X1817 => adc_samples(18179 DOWNTO 18170),
	X1818 => adc_samples(18189 DOWNTO 18180),
	X1819 => adc_samples(18199 DOWNTO 18190),
	X1820 => adc_samples(18209 DOWNTO 18200),
	X1821 => adc_samples(18219 DOWNTO 18210),
	X1822 => adc_samples(18229 DOWNTO 18220),
	X1823 => adc_samples(18239 DOWNTO 18230),
	X1824 => adc_samples(18249 DOWNTO 18240),
	X1825 => adc_samples(18259 DOWNTO 18250),
	X1826 => adc_samples(18269 DOWNTO 18260),
	X1827 => adc_samples(18279 DOWNTO 18270),
	X1828 => adc_samples(18289 DOWNTO 18280),
	X1829 => adc_samples(18299 DOWNTO 18290),
	X1830 => adc_samples(18309 DOWNTO 18300),
	X1831 => adc_samples(18319 DOWNTO 18310),
	X1832 => adc_samples(18329 DOWNTO 18320),
	X1833 => adc_samples(18339 DOWNTO 18330),
	X1834 => adc_samples(18349 DOWNTO 18340),
	X1835 => adc_samples(18359 DOWNTO 18350),
	X1836 => adc_samples(18369 DOWNTO 18360),
	X1837 => adc_samples(18379 DOWNTO 18370),
	X1838 => adc_samples(18389 DOWNTO 18380),
	X1839 => adc_samples(18399 DOWNTO 18390),
	X1840 => adc_samples(18409 DOWNTO 18400),
	X1841 => adc_samples(18419 DOWNTO 18410),
	X1842 => adc_samples(18429 DOWNTO 18420),
	X1843 => adc_samples(18439 DOWNTO 18430),
	X1844 => adc_samples(18449 DOWNTO 18440),
	X1845 => adc_samples(18459 DOWNTO 18450),
	X1846 => adc_samples(18469 DOWNTO 18460),
	X1847 => adc_samples(18479 DOWNTO 18470),
	X1848 => adc_samples(18489 DOWNTO 18480),
	X1849 => adc_samples(18499 DOWNTO 18490),
	X1850 => adc_samples(18509 DOWNTO 18500),
	X1851 => adc_samples(18519 DOWNTO 18510),
	X1852 => adc_samples(18529 DOWNTO 18520),
	X1853 => adc_samples(18539 DOWNTO 18530),
	X1854 => adc_samples(18549 DOWNTO 18540),
	X1855 => adc_samples(18559 DOWNTO 18550),
	X1856 => adc_samples(18569 DOWNTO 18560),
	X1857 => adc_samples(18579 DOWNTO 18570),
	X1858 => adc_samples(18589 DOWNTO 18580),
	X1859 => adc_samples(18599 DOWNTO 18590),
	X1860 => adc_samples(18609 DOWNTO 18600),
	X1861 => adc_samples(18619 DOWNTO 18610),
	X1862 => adc_samples(18629 DOWNTO 18620),
	X1863 => adc_samples(18639 DOWNTO 18630),
	X1864 => adc_samples(18649 DOWNTO 18640),
	X1865 => adc_samples(18659 DOWNTO 18650),
	X1866 => adc_samples(18669 DOWNTO 18660),
	X1867 => adc_samples(18679 DOWNTO 18670),
	X1868 => adc_samples(18689 DOWNTO 18680),
	X1869 => adc_samples(18699 DOWNTO 18690),
	X1870 => adc_samples(18709 DOWNTO 18700),
	X1871 => adc_samples(18719 DOWNTO 18710),
	X1872 => adc_samples(18729 DOWNTO 18720),
	X1873 => adc_samples(18739 DOWNTO 18730),
	X1874 => adc_samples(18749 DOWNTO 18740),
	X1875 => adc_samples(18759 DOWNTO 18750),
	X1876 => adc_samples(18769 DOWNTO 18760),
	X1877 => adc_samples(18779 DOWNTO 18770),
	X1878 => adc_samples(18789 DOWNTO 18780),
	X1879 => adc_samples(18799 DOWNTO 18790),
	X1880 => adc_samples(18809 DOWNTO 18800),
	X1881 => adc_samples(18819 DOWNTO 18810),
	X1882 => adc_samples(18829 DOWNTO 18820),
	X1883 => adc_samples(18839 DOWNTO 18830),
	X1884 => adc_samples(18849 DOWNTO 18840),
	X1885 => adc_samples(18859 DOWNTO 18850),
	X1886 => adc_samples(18869 DOWNTO 18860),
	X1887 => adc_samples(18879 DOWNTO 18870),
	X1888 => adc_samples(18889 DOWNTO 18880),
	X1889 => adc_samples(18899 DOWNTO 18890),
	X1890 => adc_samples(18909 DOWNTO 18900),
	X1891 => adc_samples(18919 DOWNTO 18910),
	X1892 => adc_samples(18929 DOWNTO 18920),
	X1893 => adc_samples(18939 DOWNTO 18930),
	X1894 => adc_samples(18949 DOWNTO 18940),
	X1895 => adc_samples(18959 DOWNTO 18950),
	X1896 => adc_samples(18969 DOWNTO 18960),
	X1897 => adc_samples(18979 DOWNTO 18970),
	X1898 => adc_samples(18989 DOWNTO 18980),
	X1899 => adc_samples(18999 DOWNTO 18990),
	X1900 => adc_samples(19009 DOWNTO 19000),
	X1901 => adc_samples(19019 DOWNTO 19010),
	X1902 => adc_samples(19029 DOWNTO 19020),
	X1903 => adc_samples(19039 DOWNTO 19030),
	X1904 => adc_samples(19049 DOWNTO 19040),
	X1905 => adc_samples(19059 DOWNTO 19050),
	X1906 => adc_samples(19069 DOWNTO 19060),
	X1907 => adc_samples(19079 DOWNTO 19070),
	X1908 => adc_samples(19089 DOWNTO 19080),
	X1909 => adc_samples(19099 DOWNTO 19090),
	X1910 => adc_samples(19109 DOWNTO 19100),
	X1911 => adc_samples(19119 DOWNTO 19110),
	X1912 => adc_samples(19129 DOWNTO 19120),
	X1913 => adc_samples(19139 DOWNTO 19130),
	X1914 => adc_samples(19149 DOWNTO 19140),
	X1915 => adc_samples(19159 DOWNTO 19150),
	X1916 => adc_samples(19169 DOWNTO 19160),
	X1917 => adc_samples(19179 DOWNTO 19170),
	X1918 => adc_samples(19189 DOWNTO 19180),
	X1919 => adc_samples(19199 DOWNTO 19190),
	X1920 => adc_samples(19209 DOWNTO 19200),
	X1921 => adc_samples(19219 DOWNTO 19210),
	X1922 => adc_samples(19229 DOWNTO 19220),
	X1923 => adc_samples(19239 DOWNTO 19230),
	X1924 => adc_samples(19249 DOWNTO 19240),
	X1925 => adc_samples(19259 DOWNTO 19250),
	X1926 => adc_samples(19269 DOWNTO 19260),
	X1927 => adc_samples(19279 DOWNTO 19270),
	X1928 => adc_samples(19289 DOWNTO 19280),
	X1929 => adc_samples(19299 DOWNTO 19290),
	X1930 => adc_samples(19309 DOWNTO 19300),
	X1931 => adc_samples(19319 DOWNTO 19310),
	X1932 => adc_samples(19329 DOWNTO 19320),
	X1933 => adc_samples(19339 DOWNTO 19330),
	X1934 => adc_samples(19349 DOWNTO 19340),
	X1935 => adc_samples(19359 DOWNTO 19350),
	X1936 => adc_samples(19369 DOWNTO 19360),
	X1937 => adc_samples(19379 DOWNTO 19370),
	X1938 => adc_samples(19389 DOWNTO 19380),
	X1939 => adc_samples(19399 DOWNTO 19390),
	X1940 => adc_samples(19409 DOWNTO 19400),
	X1941 => adc_samples(19419 DOWNTO 19410),
	X1942 => adc_samples(19429 DOWNTO 19420),
	X1943 => adc_samples(19439 DOWNTO 19430),
	X1944 => adc_samples(19449 DOWNTO 19440),
	X1945 => adc_samples(19459 DOWNTO 19450),
	X1946 => adc_samples(19469 DOWNTO 19460),
	X1947 => adc_samples(19479 DOWNTO 19470),
	X1948 => adc_samples(19489 DOWNTO 19480),
	X1949 => adc_samples(19499 DOWNTO 19490),
	X1950 => adc_samples(19509 DOWNTO 19500),
	X1951 => adc_samples(19519 DOWNTO 19510),
	X1952 => adc_samples(19529 DOWNTO 19520),
	X1953 => adc_samples(19539 DOWNTO 19530),
	X1954 => adc_samples(19549 DOWNTO 19540),
	X1955 => adc_samples(19559 DOWNTO 19550),
	X1956 => adc_samples(19569 DOWNTO 19560),
	X1957 => adc_samples(19579 DOWNTO 19570),
	X1958 => adc_samples(19589 DOWNTO 19580),
	X1959 => adc_samples(19599 DOWNTO 19590),
	X1960 => adc_samples(19609 DOWNTO 19600),
	X1961 => adc_samples(19619 DOWNTO 19610),
	X1962 => adc_samples(19629 DOWNTO 19620),
	X1963 => adc_samples(19639 DOWNTO 19630),
	X1964 => adc_samples(19649 DOWNTO 19640),
	X1965 => adc_samples(19659 DOWNTO 19650),
	X1966 => adc_samples(19669 DOWNTO 19660),
	X1967 => adc_samples(19679 DOWNTO 19670),
	X1968 => adc_samples(19689 DOWNTO 19680),
	X1969 => adc_samples(19699 DOWNTO 19690),
	X1970 => adc_samples(19709 DOWNTO 19700),
	X1971 => adc_samples(19719 DOWNTO 19710),
	X1972 => adc_samples(19729 DOWNTO 19720),
	X1973 => adc_samples(19739 DOWNTO 19730),
	X1974 => adc_samples(19749 DOWNTO 19740),
	X1975 => adc_samples(19759 DOWNTO 19750),
	X1976 => adc_samples(19769 DOWNTO 19760),
	X1977 => adc_samples(19779 DOWNTO 19770),
	X1978 => adc_samples(19789 DOWNTO 19780),
	X1979 => adc_samples(19799 DOWNTO 19790),
	X1980 => adc_samples(19809 DOWNTO 19800),
	X1981 => adc_samples(19819 DOWNTO 19810),
	X1982 => adc_samples(19829 DOWNTO 19820),
	X1983 => adc_samples(19839 DOWNTO 19830),
	X1984 => adc_samples(19849 DOWNTO 19840),
	X1985 => adc_samples(19859 DOWNTO 19850),
	X1986 => adc_samples(19869 DOWNTO 19860),
	X1987 => adc_samples(19879 DOWNTO 19870),
	X1988 => adc_samples(19889 DOWNTO 19880),
	X1989 => adc_samples(19899 DOWNTO 19890),
	X1990 => adc_samples(19909 DOWNTO 19900),
	X1991 => adc_samples(19919 DOWNTO 19910),
	X1992 => adc_samples(19929 DOWNTO 19920),
	X1993 => adc_samples(19939 DOWNTO 19930),
	X1994 => adc_samples(19949 DOWNTO 19940),
	X1995 => adc_samples(19959 DOWNTO 19950),
	X1996 => adc_samples(19969 DOWNTO 19960),
	X1997 => adc_samples(19979 DOWNTO 19970),
	X1998 => adc_samples(19989 DOWNTO 19980),
	X1999 => adc_samples(19999 DOWNTO 19990),
	X2000 => adc_samples(20009 DOWNTO 20000),
	X2001 => adc_samples(20019 DOWNTO 20010),
	X2002 => adc_samples(20029 DOWNTO 20020),
	X2003 => adc_samples(20039 DOWNTO 20030),
	X2004 => adc_samples(20049 DOWNTO 20040),
	X2005 => adc_samples(20059 DOWNTO 20050),
	X2006 => adc_samples(20069 DOWNTO 20060),
	X2007 => adc_samples(20079 DOWNTO 20070),
	X2008 => adc_samples(20089 DOWNTO 20080),
	X2009 => adc_samples(20099 DOWNTO 20090),
	X2010 => adc_samples(20109 DOWNTO 20100),
	X2011 => adc_samples(20119 DOWNTO 20110),
	X2012 => adc_samples(20129 DOWNTO 20120),
	X2013 => adc_samples(20139 DOWNTO 20130),
	X2014 => adc_samples(20149 DOWNTO 20140),
	X2015 => adc_samples(20159 DOWNTO 20150),
	X2016 => adc_samples(20169 DOWNTO 20160),
	X2017 => adc_samples(20179 DOWNTO 20170),
	X2018 => adc_samples(20189 DOWNTO 20180),
	X2019 => adc_samples(20199 DOWNTO 20190),
	X2020 => adc_samples(20209 DOWNTO 20200),
	X2021 => adc_samples(20219 DOWNTO 20210),
	X2022 => adc_samples(20229 DOWNTO 20220),
	X2023 => adc_samples(20239 DOWNTO 20230),
	X2024 => adc_samples(20249 DOWNTO 20240),
	X2025 => adc_samples(20259 DOWNTO 20250),
	X2026 => adc_samples(20269 DOWNTO 20260),
	X2027 => adc_samples(20279 DOWNTO 20270),
	X2028 => adc_samples(20289 DOWNTO 20280),
	X2029 => adc_samples(20299 DOWNTO 20290),
	X2030 => adc_samples(20309 DOWNTO 20300),
	X2031 => adc_samples(20319 DOWNTO 20310),
	X2032 => adc_samples(20329 DOWNTO 20320),
	X2033 => adc_samples(20339 DOWNTO 20330),
	X2034 => adc_samples(20349 DOWNTO 20340),
	X2035 => adc_samples(20359 DOWNTO 20350),
	X2036 => adc_samples(20369 DOWNTO 20360),
	X2037 => adc_samples(20379 DOWNTO 20370),
	X2038 => adc_samples(20389 DOWNTO 20380),
	X2039 => adc_samples(20399 DOWNTO 20390),
	X2040 => adc_samples(20409 DOWNTO 20400),
	X2041 => adc_samples(20419 DOWNTO 20410),
	X2042 => adc_samples(20429 DOWNTO 20420),
	X2043 => adc_samples(20439 DOWNTO 20430),
	X2044 => adc_samples(20449 DOWNTO 20440),
	X2045 => adc_samples(20459 DOWNTO 20450),
	X2046 => adc_samples(20469 DOWNTO 20460),
	X2047 => adc_samples(20479 DOWNTO 20470),
	samples_ready => samples_ready,	-- sampler has 2048 samples ready
	clk => clk,
	fft_finished => fft_finished,	-- the system is idle / can receive data
	busy => busy,	-- receiving side status
	data_ready => data_ready, -- the FFT has data ready for output / cycle data
		V0 => fft_samples(9 DOWNTO 0),
	V1 => fft_samples(19 DOWNTO 10),
	V2 => fft_samples(29 DOWNTO 20),
	V3 => fft_samples(39 DOWNTO 30),
	V4 => fft_samples(49 DOWNTO 40),
	V5 => fft_samples(59 DOWNTO 50),
	V6 => fft_samples(69 DOWNTO 60),
	V7 => fft_samples(79 DOWNTO 70),
	V8 => fft_samples(89 DOWNTO 80),
	V9 => fft_samples(99 DOWNTO 90),
	V10 => fft_samples(109 DOWNTO 100),
	V11 => fft_samples(119 DOWNTO 110),
	V12 => fft_samples(129 DOWNTO 120),
	V13 => fft_samples(139 DOWNTO 130),
	V14 => fft_samples(149 DOWNTO 140),
	V15 => fft_samples(159 DOWNTO 150)	
);

END ARCHITECTURE;