library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

ENTITY adc_sample_grabber IS
	PORT (
	ADC:    		inout std_logic_vector(11 downto 0);
	samples:   out std_logic_vector(10239 DOWNTO 0);
	clk, grab : IN std_logic;
	done : OUT STD_logic;
	sample_count : IN STD_logic_VECTOR (11 DOWNTO 0)
);
END adc_sample_grabber;

ARCHITECTURE adc_grabber OF adc_sample_grabber IS
BEGIN
	PROCESS(clk,grab,adc)
	variable temp: std_logic_vector(10239 downto 0) := (OTHERS => '0');
	BEGIN
	IF RISING_EDGE(clk) THEN
		IF (GRAB = '1') THEN
			case to_integer(unsigned(sample_count)) is
			WHEN 0 => temp(9 DOWNTO 0) := ADC(11 DOWNTO 2);
			WHEN 1 => temp(19 DOWNTO 10) := ADC(11 DOWNTO 2);
			WHEN 2 => temp(29 DOWNTO 20) := ADC(11 DOWNTO 2);
			WHEN 3 => temp(39 DOWNTO 30) := ADC(11 DOWNTO 2);
			WHEN 4 => temp(49 DOWNTO 40) := ADC(11 DOWNTO 2);
			WHEN 5 => temp(59 DOWNTO 50) := ADC(11 DOWNTO 2);
			WHEN 6 => temp(69 DOWNTO 60) := ADC(11 DOWNTO 2);
			WHEN 7 => temp(79 DOWNTO 70) := ADC(11 DOWNTO 2);
			WHEN 8 => temp(89 DOWNTO 80) := ADC(11 DOWNTO 2);
			WHEN 9 => temp(99 DOWNTO 90) := ADC(11 DOWNTO 2);
			WHEN 10 => temp(109 DOWNTO 100) := ADC(11 DOWNTO 2);
			WHEN 11 => temp(119 DOWNTO 110) := ADC(11 DOWNTO 2);
			WHEN 12 => temp(129 DOWNTO 120) := ADC(11 DOWNTO 2);
			WHEN 13 => temp(139 DOWNTO 130) := ADC(11 DOWNTO 2);
			WHEN 14 => temp(149 DOWNTO 140) := ADC(11 DOWNTO 2);
			WHEN 15 => temp(159 DOWNTO 150) := ADC(11 DOWNTO 2);
			WHEN 16 => temp(169 DOWNTO 160) := ADC(11 DOWNTO 2);
			WHEN 17 => temp(179 DOWNTO 170) := ADC(11 DOWNTO 2);
			WHEN 18 => temp(189 DOWNTO 180) := ADC(11 DOWNTO 2);
			WHEN 19 => temp(199 DOWNTO 190) := ADC(11 DOWNTO 2);
			WHEN 20 => temp(209 DOWNTO 200) := ADC(11 DOWNTO 2);
			WHEN 21 => temp(219 DOWNTO 210) := ADC(11 DOWNTO 2);
			WHEN 22 => temp(229 DOWNTO 220) := ADC(11 DOWNTO 2);
			WHEN 23 => temp(239 DOWNTO 230) := ADC(11 DOWNTO 2);
			WHEN 24 => temp(249 DOWNTO 240) := ADC(11 DOWNTO 2);
			WHEN 25 => temp(259 DOWNTO 250) := ADC(11 DOWNTO 2);
			WHEN 26 => temp(269 DOWNTO 260) := ADC(11 DOWNTO 2);
			WHEN 27 => temp(279 DOWNTO 270) := ADC(11 DOWNTO 2);
			WHEN 28 => temp(289 DOWNTO 280) := ADC(11 DOWNTO 2);
			WHEN 29 => temp(299 DOWNTO 290) := ADC(11 DOWNTO 2);
			WHEN 30 => temp(309 DOWNTO 300) := ADC(11 DOWNTO 2);
			WHEN 31 => temp(319 DOWNTO 310) := ADC(11 DOWNTO 2);
			WHEN 32 => temp(329 DOWNTO 320) := ADC(11 DOWNTO 2);
			WHEN 33 => temp(339 DOWNTO 330) := ADC(11 DOWNTO 2);
			WHEN 34 => temp(349 DOWNTO 340) := ADC(11 DOWNTO 2);
			WHEN 35 => temp(359 DOWNTO 350) := ADC(11 DOWNTO 2);
			WHEN 36 => temp(369 DOWNTO 360) := ADC(11 DOWNTO 2);
			WHEN 37 => temp(379 DOWNTO 370) := ADC(11 DOWNTO 2);
			WHEN 38 => temp(389 DOWNTO 380) := ADC(11 DOWNTO 2);
			WHEN 39 => temp(399 DOWNTO 390) := ADC(11 DOWNTO 2);
			WHEN 40 => temp(409 DOWNTO 400) := ADC(11 DOWNTO 2);
			WHEN 41 => temp(419 DOWNTO 410) := ADC(11 DOWNTO 2);
			WHEN 42 => temp(429 DOWNTO 420) := ADC(11 DOWNTO 2);
			WHEN 43 => temp(439 DOWNTO 430) := ADC(11 DOWNTO 2);
			WHEN 44 => temp(449 DOWNTO 440) := ADC(11 DOWNTO 2);
			WHEN 45 => temp(459 DOWNTO 450) := ADC(11 DOWNTO 2);
			WHEN 46 => temp(469 DOWNTO 460) := ADC(11 DOWNTO 2);
			WHEN 47 => temp(479 DOWNTO 470) := ADC(11 DOWNTO 2);
			WHEN 48 => temp(489 DOWNTO 480) := ADC(11 DOWNTO 2);
			WHEN 49 => temp(499 DOWNTO 490) := ADC(11 DOWNTO 2);
			WHEN 50 => temp(509 DOWNTO 500) := ADC(11 DOWNTO 2);
			WHEN 51 => temp(519 DOWNTO 510) := ADC(11 DOWNTO 2);
			WHEN 52 => temp(529 DOWNTO 520) := ADC(11 DOWNTO 2);
			WHEN 53 => temp(539 DOWNTO 530) := ADC(11 DOWNTO 2);
			WHEN 54 => temp(549 DOWNTO 540) := ADC(11 DOWNTO 2);
			WHEN 55 => temp(559 DOWNTO 550) := ADC(11 DOWNTO 2);
			WHEN 56 => temp(569 DOWNTO 560) := ADC(11 DOWNTO 2);
			WHEN 57 => temp(579 DOWNTO 570) := ADC(11 DOWNTO 2);
			WHEN 58 => temp(589 DOWNTO 580) := ADC(11 DOWNTO 2);
			WHEN 59 => temp(599 DOWNTO 590) := ADC(11 DOWNTO 2);
			WHEN 60 => temp(609 DOWNTO 600) := ADC(11 DOWNTO 2);
			WHEN 61 => temp(619 DOWNTO 610) := ADC(11 DOWNTO 2);
			WHEN 62 => temp(629 DOWNTO 620) := ADC(11 DOWNTO 2);
			WHEN 63 => temp(639 DOWNTO 630) := ADC(11 DOWNTO 2);
			WHEN 64 => temp(649 DOWNTO 640) := ADC(11 DOWNTO 2);
			WHEN 65 => temp(659 DOWNTO 650) := ADC(11 DOWNTO 2);
			WHEN 66 => temp(669 DOWNTO 660) := ADC(11 DOWNTO 2);
			WHEN 67 => temp(679 DOWNTO 670) := ADC(11 DOWNTO 2);
			WHEN 68 => temp(689 DOWNTO 680) := ADC(11 DOWNTO 2);
			WHEN 69 => temp(699 DOWNTO 690) := ADC(11 DOWNTO 2);
			WHEN 70 => temp(709 DOWNTO 700) := ADC(11 DOWNTO 2);
			WHEN 71 => temp(719 DOWNTO 710) := ADC(11 DOWNTO 2);
			WHEN 72 => temp(729 DOWNTO 720) := ADC(11 DOWNTO 2);
			WHEN 73 => temp(739 DOWNTO 730) := ADC(11 DOWNTO 2);
			WHEN 74 => temp(749 DOWNTO 740) := ADC(11 DOWNTO 2);
			WHEN 75 => temp(759 DOWNTO 750) := ADC(11 DOWNTO 2);
			WHEN 76 => temp(769 DOWNTO 760) := ADC(11 DOWNTO 2);
			WHEN 77 => temp(779 DOWNTO 770) := ADC(11 DOWNTO 2);
			WHEN 78 => temp(789 DOWNTO 780) := ADC(11 DOWNTO 2);
			WHEN 79 => temp(799 DOWNTO 790) := ADC(11 DOWNTO 2);
			WHEN 80 => temp(809 DOWNTO 800) := ADC(11 DOWNTO 2);
			WHEN 81 => temp(819 DOWNTO 810) := ADC(11 DOWNTO 2);
			WHEN 82 => temp(829 DOWNTO 820) := ADC(11 DOWNTO 2);
			WHEN 83 => temp(839 DOWNTO 830) := ADC(11 DOWNTO 2);
			WHEN 84 => temp(849 DOWNTO 840) := ADC(11 DOWNTO 2);
			WHEN 85 => temp(859 DOWNTO 850) := ADC(11 DOWNTO 2);
			WHEN 86 => temp(869 DOWNTO 860) := ADC(11 DOWNTO 2);
			WHEN 87 => temp(879 DOWNTO 870) := ADC(11 DOWNTO 2);
			WHEN 88 => temp(889 DOWNTO 880) := ADC(11 DOWNTO 2);
			WHEN 89 => temp(899 DOWNTO 890) := ADC(11 DOWNTO 2);
			WHEN 90 => temp(909 DOWNTO 900) := ADC(11 DOWNTO 2);
			WHEN 91 => temp(919 DOWNTO 910) := ADC(11 DOWNTO 2);
			WHEN 92 => temp(929 DOWNTO 920) := ADC(11 DOWNTO 2);
			WHEN 93 => temp(939 DOWNTO 930) := ADC(11 DOWNTO 2);
			WHEN 94 => temp(949 DOWNTO 940) := ADC(11 DOWNTO 2);
			WHEN 95 => temp(959 DOWNTO 950) := ADC(11 DOWNTO 2);
			WHEN 96 => temp(969 DOWNTO 960) := ADC(11 DOWNTO 2);
			WHEN 97 => temp(979 DOWNTO 970) := ADC(11 DOWNTO 2);
			WHEN 98 => temp(989 DOWNTO 980) := ADC(11 DOWNTO 2);
			WHEN 99 => temp(999 DOWNTO 990) := ADC(11 DOWNTO 2);
			WHEN 100 => temp(1009 DOWNTO 1000) := ADC(11 DOWNTO 2);
			WHEN 101 => temp(1019 DOWNTO 1010) := ADC(11 DOWNTO 2);
			WHEN 102 => temp(1029 DOWNTO 1020) := ADC(11 DOWNTO 2);
			WHEN 103 => temp(1039 DOWNTO 1030) := ADC(11 DOWNTO 2);
			WHEN 104 => temp(1049 DOWNTO 1040) := ADC(11 DOWNTO 2);
			WHEN 105 => temp(1059 DOWNTO 1050) := ADC(11 DOWNTO 2);
			WHEN 106 => temp(1069 DOWNTO 1060) := ADC(11 DOWNTO 2);
			WHEN 107 => temp(1079 DOWNTO 1070) := ADC(11 DOWNTO 2);
			WHEN 108 => temp(1089 DOWNTO 1080) := ADC(11 DOWNTO 2);
			WHEN 109 => temp(1099 DOWNTO 1090) := ADC(11 DOWNTO 2);
			WHEN 110 => temp(1109 DOWNTO 1100) := ADC(11 DOWNTO 2);
			WHEN 111 => temp(1119 DOWNTO 1110) := ADC(11 DOWNTO 2);
			WHEN 112 => temp(1129 DOWNTO 1120) := ADC(11 DOWNTO 2);
			WHEN 113 => temp(1139 DOWNTO 1130) := ADC(11 DOWNTO 2);
			WHEN 114 => temp(1149 DOWNTO 1140) := ADC(11 DOWNTO 2);
			WHEN 115 => temp(1159 DOWNTO 1150) := ADC(11 DOWNTO 2);
			WHEN 116 => temp(1169 DOWNTO 1160) := ADC(11 DOWNTO 2);
			WHEN 117 => temp(1179 DOWNTO 1170) := ADC(11 DOWNTO 2);
			WHEN 118 => temp(1189 DOWNTO 1180) := ADC(11 DOWNTO 2);
			WHEN 119 => temp(1199 DOWNTO 1190) := ADC(11 DOWNTO 2);
			WHEN 120 => temp(1209 DOWNTO 1200) := ADC(11 DOWNTO 2);
			WHEN 121 => temp(1219 DOWNTO 1210) := ADC(11 DOWNTO 2);
			WHEN 122 => temp(1229 DOWNTO 1220) := ADC(11 DOWNTO 2);
			WHEN 123 => temp(1239 DOWNTO 1230) := ADC(11 DOWNTO 2);
			WHEN 124 => temp(1249 DOWNTO 1240) := ADC(11 DOWNTO 2);
			WHEN 125 => temp(1259 DOWNTO 1250) := ADC(11 DOWNTO 2);
			WHEN 126 => temp(1269 DOWNTO 1260) := ADC(11 DOWNTO 2);
			WHEN 127 => temp(1279 DOWNTO 1270) := ADC(11 DOWNTO 2);
			WHEN 128 => temp(1289 DOWNTO 1280) := ADC(11 DOWNTO 2);
			WHEN 129 => temp(1299 DOWNTO 1290) := ADC(11 DOWNTO 2);
			WHEN 130 => temp(1309 DOWNTO 1300) := ADC(11 DOWNTO 2);
			WHEN 131 => temp(1319 DOWNTO 1310) := ADC(11 DOWNTO 2);
			WHEN 132 => temp(1329 DOWNTO 1320) := ADC(11 DOWNTO 2);
			WHEN 133 => temp(1339 DOWNTO 1330) := ADC(11 DOWNTO 2);
			WHEN 134 => temp(1349 DOWNTO 1340) := ADC(11 DOWNTO 2);
			WHEN 135 => temp(1359 DOWNTO 1350) := ADC(11 DOWNTO 2);
			WHEN 136 => temp(1369 DOWNTO 1360) := ADC(11 DOWNTO 2);
			WHEN 137 => temp(1379 DOWNTO 1370) := ADC(11 DOWNTO 2);
			WHEN 138 => temp(1389 DOWNTO 1380) := ADC(11 DOWNTO 2);
			WHEN 139 => temp(1399 DOWNTO 1390) := ADC(11 DOWNTO 2);
			WHEN 140 => temp(1409 DOWNTO 1400) := ADC(11 DOWNTO 2);
			WHEN 141 => temp(1419 DOWNTO 1410) := ADC(11 DOWNTO 2);
			WHEN 142 => temp(1429 DOWNTO 1420) := ADC(11 DOWNTO 2);
			WHEN 143 => temp(1439 DOWNTO 1430) := ADC(11 DOWNTO 2);
			WHEN 144 => temp(1449 DOWNTO 1440) := ADC(11 DOWNTO 2);
			WHEN 145 => temp(1459 DOWNTO 1450) := ADC(11 DOWNTO 2);
			WHEN 146 => temp(1469 DOWNTO 1460) := ADC(11 DOWNTO 2);
			WHEN 147 => temp(1479 DOWNTO 1470) := ADC(11 DOWNTO 2);
			WHEN 148 => temp(1489 DOWNTO 1480) := ADC(11 DOWNTO 2);
			WHEN 149 => temp(1499 DOWNTO 1490) := ADC(11 DOWNTO 2);
			WHEN 150 => temp(1509 DOWNTO 1500) := ADC(11 DOWNTO 2);
			WHEN 151 => temp(1519 DOWNTO 1510) := ADC(11 DOWNTO 2);
			WHEN 152 => temp(1529 DOWNTO 1520) := ADC(11 DOWNTO 2);
			WHEN 153 => temp(1539 DOWNTO 1530) := ADC(11 DOWNTO 2);
			WHEN 154 => temp(1549 DOWNTO 1540) := ADC(11 DOWNTO 2);
			WHEN 155 => temp(1559 DOWNTO 1550) := ADC(11 DOWNTO 2);
			WHEN 156 => temp(1569 DOWNTO 1560) := ADC(11 DOWNTO 2);
			WHEN 157 => temp(1579 DOWNTO 1570) := ADC(11 DOWNTO 2);
			WHEN 158 => temp(1589 DOWNTO 1580) := ADC(11 DOWNTO 2);
			WHEN 159 => temp(1599 DOWNTO 1590) := ADC(11 DOWNTO 2);
			WHEN 160 => temp(1609 DOWNTO 1600) := ADC(11 DOWNTO 2);
			WHEN 161 => temp(1619 DOWNTO 1610) := ADC(11 DOWNTO 2);
			WHEN 162 => temp(1629 DOWNTO 1620) := ADC(11 DOWNTO 2);
			WHEN 163 => temp(1639 DOWNTO 1630) := ADC(11 DOWNTO 2);
			WHEN 164 => temp(1649 DOWNTO 1640) := ADC(11 DOWNTO 2);
			WHEN 165 => temp(1659 DOWNTO 1650) := ADC(11 DOWNTO 2);
			WHEN 166 => temp(1669 DOWNTO 1660) := ADC(11 DOWNTO 2);
			WHEN 167 => temp(1679 DOWNTO 1670) := ADC(11 DOWNTO 2);
			WHEN 168 => temp(1689 DOWNTO 1680) := ADC(11 DOWNTO 2);
			WHEN 169 => temp(1699 DOWNTO 1690) := ADC(11 DOWNTO 2);
			WHEN 170 => temp(1709 DOWNTO 1700) := ADC(11 DOWNTO 2);
			WHEN 171 => temp(1719 DOWNTO 1710) := ADC(11 DOWNTO 2);
			WHEN 172 => temp(1729 DOWNTO 1720) := ADC(11 DOWNTO 2);
			WHEN 173 => temp(1739 DOWNTO 1730) := ADC(11 DOWNTO 2);
			WHEN 174 => temp(1749 DOWNTO 1740) := ADC(11 DOWNTO 2);
			WHEN 175 => temp(1759 DOWNTO 1750) := ADC(11 DOWNTO 2);
			WHEN 176 => temp(1769 DOWNTO 1760) := ADC(11 DOWNTO 2);
			WHEN 177 => temp(1779 DOWNTO 1770) := ADC(11 DOWNTO 2);
			WHEN 178 => temp(1789 DOWNTO 1780) := ADC(11 DOWNTO 2);
			WHEN 179 => temp(1799 DOWNTO 1790) := ADC(11 DOWNTO 2);
			WHEN 180 => temp(1809 DOWNTO 1800) := ADC(11 DOWNTO 2);
			WHEN 181 => temp(1819 DOWNTO 1810) := ADC(11 DOWNTO 2);
			WHEN 182 => temp(1829 DOWNTO 1820) := ADC(11 DOWNTO 2);
			WHEN 183 => temp(1839 DOWNTO 1830) := ADC(11 DOWNTO 2);
			WHEN 184 => temp(1849 DOWNTO 1840) := ADC(11 DOWNTO 2);
			WHEN 185 => temp(1859 DOWNTO 1850) := ADC(11 DOWNTO 2);
			WHEN 186 => temp(1869 DOWNTO 1860) := ADC(11 DOWNTO 2);
			WHEN 187 => temp(1879 DOWNTO 1870) := ADC(11 DOWNTO 2);
			WHEN 188 => temp(1889 DOWNTO 1880) := ADC(11 DOWNTO 2);
			WHEN 189 => temp(1899 DOWNTO 1890) := ADC(11 DOWNTO 2);
			WHEN 190 => temp(1909 DOWNTO 1900) := ADC(11 DOWNTO 2);
			WHEN 191 => temp(1919 DOWNTO 1910) := ADC(11 DOWNTO 2);
			WHEN 192 => temp(1929 DOWNTO 1920) := ADC(11 DOWNTO 2);
			WHEN 193 => temp(1939 DOWNTO 1930) := ADC(11 DOWNTO 2);
			WHEN 194 => temp(1949 DOWNTO 1940) := ADC(11 DOWNTO 2);
			WHEN 195 => temp(1959 DOWNTO 1950) := ADC(11 DOWNTO 2);
			WHEN 196 => temp(1969 DOWNTO 1960) := ADC(11 DOWNTO 2);
			WHEN 197 => temp(1979 DOWNTO 1970) := ADC(11 DOWNTO 2);
			WHEN 198 => temp(1989 DOWNTO 1980) := ADC(11 DOWNTO 2);
			WHEN 199 => temp(1999 DOWNTO 1990) := ADC(11 DOWNTO 2);
			WHEN 200 => temp(2009 DOWNTO 2000) := ADC(11 DOWNTO 2);
			WHEN 201 => temp(2019 DOWNTO 2010) := ADC(11 DOWNTO 2);
			WHEN 202 => temp(2029 DOWNTO 2020) := ADC(11 DOWNTO 2);
			WHEN 203 => temp(2039 DOWNTO 2030) := ADC(11 DOWNTO 2);
			WHEN 204 => temp(2049 DOWNTO 2040) := ADC(11 DOWNTO 2);
			WHEN 205 => temp(2059 DOWNTO 2050) := ADC(11 DOWNTO 2);
			WHEN 206 => temp(2069 DOWNTO 2060) := ADC(11 DOWNTO 2);
			WHEN 207 => temp(2079 DOWNTO 2070) := ADC(11 DOWNTO 2);
			WHEN 208 => temp(2089 DOWNTO 2080) := ADC(11 DOWNTO 2);
			WHEN 209 => temp(2099 DOWNTO 2090) := ADC(11 DOWNTO 2);
			WHEN 210 => temp(2109 DOWNTO 2100) := ADC(11 DOWNTO 2);
			WHEN 211 => temp(2119 DOWNTO 2110) := ADC(11 DOWNTO 2);
			WHEN 212 => temp(2129 DOWNTO 2120) := ADC(11 DOWNTO 2);
			WHEN 213 => temp(2139 DOWNTO 2130) := ADC(11 DOWNTO 2);
			WHEN 214 => temp(2149 DOWNTO 2140) := ADC(11 DOWNTO 2);
			WHEN 215 => temp(2159 DOWNTO 2150) := ADC(11 DOWNTO 2);
			WHEN 216 => temp(2169 DOWNTO 2160) := ADC(11 DOWNTO 2);
			WHEN 217 => temp(2179 DOWNTO 2170) := ADC(11 DOWNTO 2);
			WHEN 218 => temp(2189 DOWNTO 2180) := ADC(11 DOWNTO 2);
			WHEN 219 => temp(2199 DOWNTO 2190) := ADC(11 DOWNTO 2);
			WHEN 220 => temp(2209 DOWNTO 2200) := ADC(11 DOWNTO 2);
			WHEN 221 => temp(2219 DOWNTO 2210) := ADC(11 DOWNTO 2);
			WHEN 222 => temp(2229 DOWNTO 2220) := ADC(11 DOWNTO 2);
			WHEN 223 => temp(2239 DOWNTO 2230) := ADC(11 DOWNTO 2);
			WHEN 224 => temp(2249 DOWNTO 2240) := ADC(11 DOWNTO 2);
			WHEN 225 => temp(2259 DOWNTO 2250) := ADC(11 DOWNTO 2);
			WHEN 226 => temp(2269 DOWNTO 2260) := ADC(11 DOWNTO 2);
			WHEN 227 => temp(2279 DOWNTO 2270) := ADC(11 DOWNTO 2);
			WHEN 228 => temp(2289 DOWNTO 2280) := ADC(11 DOWNTO 2);
			WHEN 229 => temp(2299 DOWNTO 2290) := ADC(11 DOWNTO 2);
			WHEN 230 => temp(2309 DOWNTO 2300) := ADC(11 DOWNTO 2);
			WHEN 231 => temp(2319 DOWNTO 2310) := ADC(11 DOWNTO 2);
			WHEN 232 => temp(2329 DOWNTO 2320) := ADC(11 DOWNTO 2);
			WHEN 233 => temp(2339 DOWNTO 2330) := ADC(11 DOWNTO 2);
			WHEN 234 => temp(2349 DOWNTO 2340) := ADC(11 DOWNTO 2);
			WHEN 235 => temp(2359 DOWNTO 2350) := ADC(11 DOWNTO 2);
			WHEN 236 => temp(2369 DOWNTO 2360) := ADC(11 DOWNTO 2);
			WHEN 237 => temp(2379 DOWNTO 2370) := ADC(11 DOWNTO 2);
			WHEN 238 => temp(2389 DOWNTO 2380) := ADC(11 DOWNTO 2);
			WHEN 239 => temp(2399 DOWNTO 2390) := ADC(11 DOWNTO 2);
			WHEN 240 => temp(2409 DOWNTO 2400) := ADC(11 DOWNTO 2);
			WHEN 241 => temp(2419 DOWNTO 2410) := ADC(11 DOWNTO 2);
			WHEN 242 => temp(2429 DOWNTO 2420) := ADC(11 DOWNTO 2);
			WHEN 243 => temp(2439 DOWNTO 2430) := ADC(11 DOWNTO 2);
			WHEN 244 => temp(2449 DOWNTO 2440) := ADC(11 DOWNTO 2);
			WHEN 245 => temp(2459 DOWNTO 2450) := ADC(11 DOWNTO 2);
			WHEN 246 => temp(2469 DOWNTO 2460) := ADC(11 DOWNTO 2);
			WHEN 247 => temp(2479 DOWNTO 2470) := ADC(11 DOWNTO 2);
			WHEN 248 => temp(2489 DOWNTO 2480) := ADC(11 DOWNTO 2);
			WHEN 249 => temp(2499 DOWNTO 2490) := ADC(11 DOWNTO 2);
			WHEN 250 => temp(2509 DOWNTO 2500) := ADC(11 DOWNTO 2);
			WHEN 251 => temp(2519 DOWNTO 2510) := ADC(11 DOWNTO 2);
			WHEN 252 => temp(2529 DOWNTO 2520) := ADC(11 DOWNTO 2);
			WHEN 253 => temp(2539 DOWNTO 2530) := ADC(11 DOWNTO 2);
			WHEN 254 => temp(2549 DOWNTO 2540) := ADC(11 DOWNTO 2);
			WHEN 255 => temp(2559 DOWNTO 2550) := ADC(11 DOWNTO 2);
			WHEN 256 => temp(2569 DOWNTO 2560) := ADC(11 DOWNTO 2);
			WHEN 257 => temp(2579 DOWNTO 2570) := ADC(11 DOWNTO 2);
			WHEN 258 => temp(2589 DOWNTO 2580) := ADC(11 DOWNTO 2);
			WHEN 259 => temp(2599 DOWNTO 2590) := ADC(11 DOWNTO 2);
			WHEN 260 => temp(2609 DOWNTO 2600) := ADC(11 DOWNTO 2);
			WHEN 261 => temp(2619 DOWNTO 2610) := ADC(11 DOWNTO 2);
			WHEN 262 => temp(2629 DOWNTO 2620) := ADC(11 DOWNTO 2);
			WHEN 263 => temp(2639 DOWNTO 2630) := ADC(11 DOWNTO 2);
			WHEN 264 => temp(2649 DOWNTO 2640) := ADC(11 DOWNTO 2);
			WHEN 265 => temp(2659 DOWNTO 2650) := ADC(11 DOWNTO 2);
			WHEN 266 => temp(2669 DOWNTO 2660) := ADC(11 DOWNTO 2);
			WHEN 267 => temp(2679 DOWNTO 2670) := ADC(11 DOWNTO 2);
			WHEN 268 => temp(2689 DOWNTO 2680) := ADC(11 DOWNTO 2);
			WHEN 269 => temp(2699 DOWNTO 2690) := ADC(11 DOWNTO 2);
			WHEN 270 => temp(2709 DOWNTO 2700) := ADC(11 DOWNTO 2);
			WHEN 271 => temp(2719 DOWNTO 2710) := ADC(11 DOWNTO 2);
			WHEN 272 => temp(2729 DOWNTO 2720) := ADC(11 DOWNTO 2);
			WHEN 273 => temp(2739 DOWNTO 2730) := ADC(11 DOWNTO 2);
			WHEN 274 => temp(2749 DOWNTO 2740) := ADC(11 DOWNTO 2);
			WHEN 275 => temp(2759 DOWNTO 2750) := ADC(11 DOWNTO 2);
			WHEN 276 => temp(2769 DOWNTO 2760) := ADC(11 DOWNTO 2);
			WHEN 277 => temp(2779 DOWNTO 2770) := ADC(11 DOWNTO 2);
			WHEN 278 => temp(2789 DOWNTO 2780) := ADC(11 DOWNTO 2);
			WHEN 279 => temp(2799 DOWNTO 2790) := ADC(11 DOWNTO 2);
			WHEN 280 => temp(2809 DOWNTO 2800) := ADC(11 DOWNTO 2);
			WHEN 281 => temp(2819 DOWNTO 2810) := ADC(11 DOWNTO 2);
			WHEN 282 => temp(2829 DOWNTO 2820) := ADC(11 DOWNTO 2);
			WHEN 283 => temp(2839 DOWNTO 2830) := ADC(11 DOWNTO 2);
			WHEN 284 => temp(2849 DOWNTO 2840) := ADC(11 DOWNTO 2);
			WHEN 285 => temp(2859 DOWNTO 2850) := ADC(11 DOWNTO 2);
			WHEN 286 => temp(2869 DOWNTO 2860) := ADC(11 DOWNTO 2);
			WHEN 287 => temp(2879 DOWNTO 2870) := ADC(11 DOWNTO 2);
			WHEN 288 => temp(2889 DOWNTO 2880) := ADC(11 DOWNTO 2);
			WHEN 289 => temp(2899 DOWNTO 2890) := ADC(11 DOWNTO 2);
			WHEN 290 => temp(2909 DOWNTO 2900) := ADC(11 DOWNTO 2);
			WHEN 291 => temp(2919 DOWNTO 2910) := ADC(11 DOWNTO 2);
			WHEN 292 => temp(2929 DOWNTO 2920) := ADC(11 DOWNTO 2);
			WHEN 293 => temp(2939 DOWNTO 2930) := ADC(11 DOWNTO 2);
			WHEN 294 => temp(2949 DOWNTO 2940) := ADC(11 DOWNTO 2);
			WHEN 295 => temp(2959 DOWNTO 2950) := ADC(11 DOWNTO 2);
			WHEN 296 => temp(2969 DOWNTO 2960) := ADC(11 DOWNTO 2);
			WHEN 297 => temp(2979 DOWNTO 2970) := ADC(11 DOWNTO 2);
			WHEN 298 => temp(2989 DOWNTO 2980) := ADC(11 DOWNTO 2);
			WHEN 299 => temp(2999 DOWNTO 2990) := ADC(11 DOWNTO 2);
			WHEN 300 => temp(3009 DOWNTO 3000) := ADC(11 DOWNTO 2);
			WHEN 301 => temp(3019 DOWNTO 3010) := ADC(11 DOWNTO 2);
			WHEN 302 => temp(3029 DOWNTO 3020) := ADC(11 DOWNTO 2);
			WHEN 303 => temp(3039 DOWNTO 3030) := ADC(11 DOWNTO 2);
			WHEN 304 => temp(3049 DOWNTO 3040) := ADC(11 DOWNTO 2);
			WHEN 305 => temp(3059 DOWNTO 3050) := ADC(11 DOWNTO 2);
			WHEN 306 => temp(3069 DOWNTO 3060) := ADC(11 DOWNTO 2);
			WHEN 307 => temp(3079 DOWNTO 3070) := ADC(11 DOWNTO 2);
			WHEN 308 => temp(3089 DOWNTO 3080) := ADC(11 DOWNTO 2);
			WHEN 309 => temp(3099 DOWNTO 3090) := ADC(11 DOWNTO 2);
			WHEN 310 => temp(3109 DOWNTO 3100) := ADC(11 DOWNTO 2);
			WHEN 311 => temp(3119 DOWNTO 3110) := ADC(11 DOWNTO 2);
			WHEN 312 => temp(3129 DOWNTO 3120) := ADC(11 DOWNTO 2);
			WHEN 313 => temp(3139 DOWNTO 3130) := ADC(11 DOWNTO 2);
			WHEN 314 => temp(3149 DOWNTO 3140) := ADC(11 DOWNTO 2);
			WHEN 315 => temp(3159 DOWNTO 3150) := ADC(11 DOWNTO 2);
			WHEN 316 => temp(3169 DOWNTO 3160) := ADC(11 DOWNTO 2);
			WHEN 317 => temp(3179 DOWNTO 3170) := ADC(11 DOWNTO 2);
			WHEN 318 => temp(3189 DOWNTO 3180) := ADC(11 DOWNTO 2);
			WHEN 319 => temp(3199 DOWNTO 3190) := ADC(11 DOWNTO 2);
			WHEN 320 => temp(3209 DOWNTO 3200) := ADC(11 DOWNTO 2);
			WHEN 321 => temp(3219 DOWNTO 3210) := ADC(11 DOWNTO 2);
			WHEN 322 => temp(3229 DOWNTO 3220) := ADC(11 DOWNTO 2);
			WHEN 323 => temp(3239 DOWNTO 3230) := ADC(11 DOWNTO 2);
			WHEN 324 => temp(3249 DOWNTO 3240) := ADC(11 DOWNTO 2);
			WHEN 325 => temp(3259 DOWNTO 3250) := ADC(11 DOWNTO 2);
			WHEN 326 => temp(3269 DOWNTO 3260) := ADC(11 DOWNTO 2);
			WHEN 327 => temp(3279 DOWNTO 3270) := ADC(11 DOWNTO 2);
			WHEN 328 => temp(3289 DOWNTO 3280) := ADC(11 DOWNTO 2);
			WHEN 329 => temp(3299 DOWNTO 3290) := ADC(11 DOWNTO 2);
			WHEN 330 => temp(3309 DOWNTO 3300) := ADC(11 DOWNTO 2);
			WHEN 331 => temp(3319 DOWNTO 3310) := ADC(11 DOWNTO 2);
			WHEN 332 => temp(3329 DOWNTO 3320) := ADC(11 DOWNTO 2);
			WHEN 333 => temp(3339 DOWNTO 3330) := ADC(11 DOWNTO 2);
			WHEN 334 => temp(3349 DOWNTO 3340) := ADC(11 DOWNTO 2);
			WHEN 335 => temp(3359 DOWNTO 3350) := ADC(11 DOWNTO 2);
			WHEN 336 => temp(3369 DOWNTO 3360) := ADC(11 DOWNTO 2);
			WHEN 337 => temp(3379 DOWNTO 3370) := ADC(11 DOWNTO 2);
			WHEN 338 => temp(3389 DOWNTO 3380) := ADC(11 DOWNTO 2);
			WHEN 339 => temp(3399 DOWNTO 3390) := ADC(11 DOWNTO 2);
			WHEN 340 => temp(3409 DOWNTO 3400) := ADC(11 DOWNTO 2);
			WHEN 341 => temp(3419 DOWNTO 3410) := ADC(11 DOWNTO 2);
			WHEN 342 => temp(3429 DOWNTO 3420) := ADC(11 DOWNTO 2);
			WHEN 343 => temp(3439 DOWNTO 3430) := ADC(11 DOWNTO 2);
			WHEN 344 => temp(3449 DOWNTO 3440) := ADC(11 DOWNTO 2);
			WHEN 345 => temp(3459 DOWNTO 3450) := ADC(11 DOWNTO 2);
			WHEN 346 => temp(3469 DOWNTO 3460) := ADC(11 DOWNTO 2);
			WHEN 347 => temp(3479 DOWNTO 3470) := ADC(11 DOWNTO 2);
			WHEN 348 => temp(3489 DOWNTO 3480) := ADC(11 DOWNTO 2);
			WHEN 349 => temp(3499 DOWNTO 3490) := ADC(11 DOWNTO 2);
			WHEN 350 => temp(3509 DOWNTO 3500) := ADC(11 DOWNTO 2);
			WHEN 351 => temp(3519 DOWNTO 3510) := ADC(11 DOWNTO 2);
			WHEN 352 => temp(3529 DOWNTO 3520) := ADC(11 DOWNTO 2);
			WHEN 353 => temp(3539 DOWNTO 3530) := ADC(11 DOWNTO 2);
			WHEN 354 => temp(3549 DOWNTO 3540) := ADC(11 DOWNTO 2);
			WHEN 355 => temp(3559 DOWNTO 3550) := ADC(11 DOWNTO 2);
			WHEN 356 => temp(3569 DOWNTO 3560) := ADC(11 DOWNTO 2);
			WHEN 357 => temp(3579 DOWNTO 3570) := ADC(11 DOWNTO 2);
			WHEN 358 => temp(3589 DOWNTO 3580) := ADC(11 DOWNTO 2);
			WHEN 359 => temp(3599 DOWNTO 3590) := ADC(11 DOWNTO 2);
			WHEN 360 => temp(3609 DOWNTO 3600) := ADC(11 DOWNTO 2);
			WHEN 361 => temp(3619 DOWNTO 3610) := ADC(11 DOWNTO 2);
			WHEN 362 => temp(3629 DOWNTO 3620) := ADC(11 DOWNTO 2);
			WHEN 363 => temp(3639 DOWNTO 3630) := ADC(11 DOWNTO 2);
			WHEN 364 => temp(3649 DOWNTO 3640) := ADC(11 DOWNTO 2);
			WHEN 365 => temp(3659 DOWNTO 3650) := ADC(11 DOWNTO 2);
			WHEN 366 => temp(3669 DOWNTO 3660) := ADC(11 DOWNTO 2);
			WHEN 367 => temp(3679 DOWNTO 3670) := ADC(11 DOWNTO 2);
			WHEN 368 => temp(3689 DOWNTO 3680) := ADC(11 DOWNTO 2);
			WHEN 369 => temp(3699 DOWNTO 3690) := ADC(11 DOWNTO 2);
			WHEN 370 => temp(3709 DOWNTO 3700) := ADC(11 DOWNTO 2);
			WHEN 371 => temp(3719 DOWNTO 3710) := ADC(11 DOWNTO 2);
			WHEN 372 => temp(3729 DOWNTO 3720) := ADC(11 DOWNTO 2);
			WHEN 373 => temp(3739 DOWNTO 3730) := ADC(11 DOWNTO 2);
			WHEN 374 => temp(3749 DOWNTO 3740) := ADC(11 DOWNTO 2);
			WHEN 375 => temp(3759 DOWNTO 3750) := ADC(11 DOWNTO 2);
			WHEN 376 => temp(3769 DOWNTO 3760) := ADC(11 DOWNTO 2);
			WHEN 377 => temp(3779 DOWNTO 3770) := ADC(11 DOWNTO 2);
			WHEN 378 => temp(3789 DOWNTO 3780) := ADC(11 DOWNTO 2);
			WHEN 379 => temp(3799 DOWNTO 3790) := ADC(11 DOWNTO 2);
			WHEN 380 => temp(3809 DOWNTO 3800) := ADC(11 DOWNTO 2);
			WHEN 381 => temp(3819 DOWNTO 3810) := ADC(11 DOWNTO 2);
			WHEN 382 => temp(3829 DOWNTO 3820) := ADC(11 DOWNTO 2);
			WHEN 383 => temp(3839 DOWNTO 3830) := ADC(11 DOWNTO 2);
			WHEN 384 => temp(3849 DOWNTO 3840) := ADC(11 DOWNTO 2);
			WHEN 385 => temp(3859 DOWNTO 3850) := ADC(11 DOWNTO 2);
			WHEN 386 => temp(3869 DOWNTO 3860) := ADC(11 DOWNTO 2);
			WHEN 387 => temp(3879 DOWNTO 3870) := ADC(11 DOWNTO 2);
			WHEN 388 => temp(3889 DOWNTO 3880) := ADC(11 DOWNTO 2);
			WHEN 389 => temp(3899 DOWNTO 3890) := ADC(11 DOWNTO 2);
			WHEN 390 => temp(3909 DOWNTO 3900) := ADC(11 DOWNTO 2);
			WHEN 391 => temp(3919 DOWNTO 3910) := ADC(11 DOWNTO 2);
			WHEN 392 => temp(3929 DOWNTO 3920) := ADC(11 DOWNTO 2);
			WHEN 393 => temp(3939 DOWNTO 3930) := ADC(11 DOWNTO 2);
			WHEN 394 => temp(3949 DOWNTO 3940) := ADC(11 DOWNTO 2);
			WHEN 395 => temp(3959 DOWNTO 3950) := ADC(11 DOWNTO 2);
			WHEN 396 => temp(3969 DOWNTO 3960) := ADC(11 DOWNTO 2);
			WHEN 397 => temp(3979 DOWNTO 3970) := ADC(11 DOWNTO 2);
			WHEN 398 => temp(3989 DOWNTO 3980) := ADC(11 DOWNTO 2);
			WHEN 399 => temp(3999 DOWNTO 3990) := ADC(11 DOWNTO 2);
			WHEN 400 => temp(4009 DOWNTO 4000) := ADC(11 DOWNTO 2);
			WHEN 401 => temp(4019 DOWNTO 4010) := ADC(11 DOWNTO 2);
			WHEN 402 => temp(4029 DOWNTO 4020) := ADC(11 DOWNTO 2);
			WHEN 403 => temp(4039 DOWNTO 4030) := ADC(11 DOWNTO 2);
			WHEN 404 => temp(4049 DOWNTO 4040) := ADC(11 DOWNTO 2);
			WHEN 405 => temp(4059 DOWNTO 4050) := ADC(11 DOWNTO 2);
			WHEN 406 => temp(4069 DOWNTO 4060) := ADC(11 DOWNTO 2);
			WHEN 407 => temp(4079 DOWNTO 4070) := ADC(11 DOWNTO 2);
			WHEN 408 => temp(4089 DOWNTO 4080) := ADC(11 DOWNTO 2);
			WHEN 409 => temp(4099 DOWNTO 4090) := ADC(11 DOWNTO 2);
			WHEN 410 => temp(4109 DOWNTO 4100) := ADC(11 DOWNTO 2);
			WHEN 411 => temp(4119 DOWNTO 4110) := ADC(11 DOWNTO 2);
			WHEN 412 => temp(4129 DOWNTO 4120) := ADC(11 DOWNTO 2);
			WHEN 413 => temp(4139 DOWNTO 4130) := ADC(11 DOWNTO 2);
			WHEN 414 => temp(4149 DOWNTO 4140) := ADC(11 DOWNTO 2);
			WHEN 415 => temp(4159 DOWNTO 4150) := ADC(11 DOWNTO 2);
			WHEN 416 => temp(4169 DOWNTO 4160) := ADC(11 DOWNTO 2);
			WHEN 417 => temp(4179 DOWNTO 4170) := ADC(11 DOWNTO 2);
			WHEN 418 => temp(4189 DOWNTO 4180) := ADC(11 DOWNTO 2);
			WHEN 419 => temp(4199 DOWNTO 4190) := ADC(11 DOWNTO 2);
			WHEN 420 => temp(4209 DOWNTO 4200) := ADC(11 DOWNTO 2);
			WHEN 421 => temp(4219 DOWNTO 4210) := ADC(11 DOWNTO 2);
			WHEN 422 => temp(4229 DOWNTO 4220) := ADC(11 DOWNTO 2);
			WHEN 423 => temp(4239 DOWNTO 4230) := ADC(11 DOWNTO 2);
			WHEN 424 => temp(4249 DOWNTO 4240) := ADC(11 DOWNTO 2);
			WHEN 425 => temp(4259 DOWNTO 4250) := ADC(11 DOWNTO 2);
			WHEN 426 => temp(4269 DOWNTO 4260) := ADC(11 DOWNTO 2);
			WHEN 427 => temp(4279 DOWNTO 4270) := ADC(11 DOWNTO 2);
			WHEN 428 => temp(4289 DOWNTO 4280) := ADC(11 DOWNTO 2);
			WHEN 429 => temp(4299 DOWNTO 4290) := ADC(11 DOWNTO 2);
			WHEN 430 => temp(4309 DOWNTO 4300) := ADC(11 DOWNTO 2);
			WHEN 431 => temp(4319 DOWNTO 4310) := ADC(11 DOWNTO 2);
			WHEN 432 => temp(4329 DOWNTO 4320) := ADC(11 DOWNTO 2);
			WHEN 433 => temp(4339 DOWNTO 4330) := ADC(11 DOWNTO 2);
			WHEN 434 => temp(4349 DOWNTO 4340) := ADC(11 DOWNTO 2);
			WHEN 435 => temp(4359 DOWNTO 4350) := ADC(11 DOWNTO 2);
			WHEN 436 => temp(4369 DOWNTO 4360) := ADC(11 DOWNTO 2);
			WHEN 437 => temp(4379 DOWNTO 4370) := ADC(11 DOWNTO 2);
			WHEN 438 => temp(4389 DOWNTO 4380) := ADC(11 DOWNTO 2);
			WHEN 439 => temp(4399 DOWNTO 4390) := ADC(11 DOWNTO 2);
			WHEN 440 => temp(4409 DOWNTO 4400) := ADC(11 DOWNTO 2);
			WHEN 441 => temp(4419 DOWNTO 4410) := ADC(11 DOWNTO 2);
			WHEN 442 => temp(4429 DOWNTO 4420) := ADC(11 DOWNTO 2);
			WHEN 443 => temp(4439 DOWNTO 4430) := ADC(11 DOWNTO 2);
			WHEN 444 => temp(4449 DOWNTO 4440) := ADC(11 DOWNTO 2);
			WHEN 445 => temp(4459 DOWNTO 4450) := ADC(11 DOWNTO 2);
			WHEN 446 => temp(4469 DOWNTO 4460) := ADC(11 DOWNTO 2);
			WHEN 447 => temp(4479 DOWNTO 4470) := ADC(11 DOWNTO 2);
			WHEN 448 => temp(4489 DOWNTO 4480) := ADC(11 DOWNTO 2);
			WHEN 449 => temp(4499 DOWNTO 4490) := ADC(11 DOWNTO 2);
			WHEN 450 => temp(4509 DOWNTO 4500) := ADC(11 DOWNTO 2);
			WHEN 451 => temp(4519 DOWNTO 4510) := ADC(11 DOWNTO 2);
			WHEN 452 => temp(4529 DOWNTO 4520) := ADC(11 DOWNTO 2);
			WHEN 453 => temp(4539 DOWNTO 4530) := ADC(11 DOWNTO 2);
			WHEN 454 => temp(4549 DOWNTO 4540) := ADC(11 DOWNTO 2);
			WHEN 455 => temp(4559 DOWNTO 4550) := ADC(11 DOWNTO 2);
			WHEN 456 => temp(4569 DOWNTO 4560) := ADC(11 DOWNTO 2);
			WHEN 457 => temp(4579 DOWNTO 4570) := ADC(11 DOWNTO 2);
			WHEN 458 => temp(4589 DOWNTO 4580) := ADC(11 DOWNTO 2);
			WHEN 459 => temp(4599 DOWNTO 4590) := ADC(11 DOWNTO 2);
			WHEN 460 => temp(4609 DOWNTO 4600) := ADC(11 DOWNTO 2);
			WHEN 461 => temp(4619 DOWNTO 4610) := ADC(11 DOWNTO 2);
			WHEN 462 => temp(4629 DOWNTO 4620) := ADC(11 DOWNTO 2);
			WHEN 463 => temp(4639 DOWNTO 4630) := ADC(11 DOWNTO 2);
			WHEN 464 => temp(4649 DOWNTO 4640) := ADC(11 DOWNTO 2);
			WHEN 465 => temp(4659 DOWNTO 4650) := ADC(11 DOWNTO 2);
			WHEN 466 => temp(4669 DOWNTO 4660) := ADC(11 DOWNTO 2);
			WHEN 467 => temp(4679 DOWNTO 4670) := ADC(11 DOWNTO 2);
			WHEN 468 => temp(4689 DOWNTO 4680) := ADC(11 DOWNTO 2);
			WHEN 469 => temp(4699 DOWNTO 4690) := ADC(11 DOWNTO 2);
			WHEN 470 => temp(4709 DOWNTO 4700) := ADC(11 DOWNTO 2);
			WHEN 471 => temp(4719 DOWNTO 4710) := ADC(11 DOWNTO 2);
			WHEN 472 => temp(4729 DOWNTO 4720) := ADC(11 DOWNTO 2);
			WHEN 473 => temp(4739 DOWNTO 4730) := ADC(11 DOWNTO 2);
			WHEN 474 => temp(4749 DOWNTO 4740) := ADC(11 DOWNTO 2);
			WHEN 475 => temp(4759 DOWNTO 4750) := ADC(11 DOWNTO 2);
			WHEN 476 => temp(4769 DOWNTO 4760) := ADC(11 DOWNTO 2);
			WHEN 477 => temp(4779 DOWNTO 4770) := ADC(11 DOWNTO 2);
			WHEN 478 => temp(4789 DOWNTO 4780) := ADC(11 DOWNTO 2);
			WHEN 479 => temp(4799 DOWNTO 4790) := ADC(11 DOWNTO 2);
			WHEN 480 => temp(4809 DOWNTO 4800) := ADC(11 DOWNTO 2);
			WHEN 481 => temp(4819 DOWNTO 4810) := ADC(11 DOWNTO 2);
			WHEN 482 => temp(4829 DOWNTO 4820) := ADC(11 DOWNTO 2);
			WHEN 483 => temp(4839 DOWNTO 4830) := ADC(11 DOWNTO 2);
			WHEN 484 => temp(4849 DOWNTO 4840) := ADC(11 DOWNTO 2);
			WHEN 485 => temp(4859 DOWNTO 4850) := ADC(11 DOWNTO 2);
			WHEN 486 => temp(4869 DOWNTO 4860) := ADC(11 DOWNTO 2);
			WHEN 487 => temp(4879 DOWNTO 4870) := ADC(11 DOWNTO 2);
			WHEN 488 => temp(4889 DOWNTO 4880) := ADC(11 DOWNTO 2);
			WHEN 489 => temp(4899 DOWNTO 4890) := ADC(11 DOWNTO 2);
			WHEN 490 => temp(4909 DOWNTO 4900) := ADC(11 DOWNTO 2);
			WHEN 491 => temp(4919 DOWNTO 4910) := ADC(11 DOWNTO 2);
			WHEN 492 => temp(4929 DOWNTO 4920) := ADC(11 DOWNTO 2);
			WHEN 493 => temp(4939 DOWNTO 4930) := ADC(11 DOWNTO 2);
			WHEN 494 => temp(4949 DOWNTO 4940) := ADC(11 DOWNTO 2);
			WHEN 495 => temp(4959 DOWNTO 4950) := ADC(11 DOWNTO 2);
			WHEN 496 => temp(4969 DOWNTO 4960) := ADC(11 DOWNTO 2);
			WHEN 497 => temp(4979 DOWNTO 4970) := ADC(11 DOWNTO 2);
			WHEN 498 => temp(4989 DOWNTO 4980) := ADC(11 DOWNTO 2);
			WHEN 499 => temp(4999 DOWNTO 4990) := ADC(11 DOWNTO 2);
			WHEN 500 => temp(5009 DOWNTO 5000) := ADC(11 DOWNTO 2);
			WHEN 501 => temp(5019 DOWNTO 5010) := ADC(11 DOWNTO 2);
			WHEN 502 => temp(5029 DOWNTO 5020) := ADC(11 DOWNTO 2);
			WHEN 503 => temp(5039 DOWNTO 5030) := ADC(11 DOWNTO 2);
			WHEN 504 => temp(5049 DOWNTO 5040) := ADC(11 DOWNTO 2);
			WHEN 505 => temp(5059 DOWNTO 5050) := ADC(11 DOWNTO 2);
			WHEN 506 => temp(5069 DOWNTO 5060) := ADC(11 DOWNTO 2);
			WHEN 507 => temp(5079 DOWNTO 5070) := ADC(11 DOWNTO 2);
			WHEN 508 => temp(5089 DOWNTO 5080) := ADC(11 DOWNTO 2);
			WHEN 509 => temp(5099 DOWNTO 5090) := ADC(11 DOWNTO 2);
			WHEN 510 => temp(5109 DOWNTO 5100) := ADC(11 DOWNTO 2);
			WHEN 511 => temp(5119 DOWNTO 5110) := ADC(11 DOWNTO 2);
			WHEN 512 => temp(5129 DOWNTO 5120) := ADC(11 DOWNTO 2);
			WHEN 513 => temp(5139 DOWNTO 5130) := ADC(11 DOWNTO 2);
			WHEN 514 => temp(5149 DOWNTO 5140) := ADC(11 DOWNTO 2);
			WHEN 515 => temp(5159 DOWNTO 5150) := ADC(11 DOWNTO 2);
			WHEN 516 => temp(5169 DOWNTO 5160) := ADC(11 DOWNTO 2);
			WHEN 517 => temp(5179 DOWNTO 5170) := ADC(11 DOWNTO 2);
			WHEN 518 => temp(5189 DOWNTO 5180) := ADC(11 DOWNTO 2);
			WHEN 519 => temp(5199 DOWNTO 5190) := ADC(11 DOWNTO 2);
			WHEN 520 => temp(5209 DOWNTO 5200) := ADC(11 DOWNTO 2);
			WHEN 521 => temp(5219 DOWNTO 5210) := ADC(11 DOWNTO 2);
			WHEN 522 => temp(5229 DOWNTO 5220) := ADC(11 DOWNTO 2);
			WHEN 523 => temp(5239 DOWNTO 5230) := ADC(11 DOWNTO 2);
			WHEN 524 => temp(5249 DOWNTO 5240) := ADC(11 DOWNTO 2);
			WHEN 525 => temp(5259 DOWNTO 5250) := ADC(11 DOWNTO 2);
			WHEN 526 => temp(5269 DOWNTO 5260) := ADC(11 DOWNTO 2);
			WHEN 527 => temp(5279 DOWNTO 5270) := ADC(11 DOWNTO 2);
			WHEN 528 => temp(5289 DOWNTO 5280) := ADC(11 DOWNTO 2);
			WHEN 529 => temp(5299 DOWNTO 5290) := ADC(11 DOWNTO 2);
			WHEN 530 => temp(5309 DOWNTO 5300) := ADC(11 DOWNTO 2);
			WHEN 531 => temp(5319 DOWNTO 5310) := ADC(11 DOWNTO 2);
			WHEN 532 => temp(5329 DOWNTO 5320) := ADC(11 DOWNTO 2);
			WHEN 533 => temp(5339 DOWNTO 5330) := ADC(11 DOWNTO 2);
			WHEN 534 => temp(5349 DOWNTO 5340) := ADC(11 DOWNTO 2);
			WHEN 535 => temp(5359 DOWNTO 5350) := ADC(11 DOWNTO 2);
			WHEN 536 => temp(5369 DOWNTO 5360) := ADC(11 DOWNTO 2);
			WHEN 537 => temp(5379 DOWNTO 5370) := ADC(11 DOWNTO 2);
			WHEN 538 => temp(5389 DOWNTO 5380) := ADC(11 DOWNTO 2);
			WHEN 539 => temp(5399 DOWNTO 5390) := ADC(11 DOWNTO 2);
			WHEN 540 => temp(5409 DOWNTO 5400) := ADC(11 DOWNTO 2);
			WHEN 541 => temp(5419 DOWNTO 5410) := ADC(11 DOWNTO 2);
			WHEN 542 => temp(5429 DOWNTO 5420) := ADC(11 DOWNTO 2);
			WHEN 543 => temp(5439 DOWNTO 5430) := ADC(11 DOWNTO 2);
			WHEN 544 => temp(5449 DOWNTO 5440) := ADC(11 DOWNTO 2);
			WHEN 545 => temp(5459 DOWNTO 5450) := ADC(11 DOWNTO 2);
			WHEN 546 => temp(5469 DOWNTO 5460) := ADC(11 DOWNTO 2);
			WHEN 547 => temp(5479 DOWNTO 5470) := ADC(11 DOWNTO 2);
			WHEN 548 => temp(5489 DOWNTO 5480) := ADC(11 DOWNTO 2);
			WHEN 549 => temp(5499 DOWNTO 5490) := ADC(11 DOWNTO 2);
			WHEN 550 => temp(5509 DOWNTO 5500) := ADC(11 DOWNTO 2);
			WHEN 551 => temp(5519 DOWNTO 5510) := ADC(11 DOWNTO 2);
			WHEN 552 => temp(5529 DOWNTO 5520) := ADC(11 DOWNTO 2);
			WHEN 553 => temp(5539 DOWNTO 5530) := ADC(11 DOWNTO 2);
			WHEN 554 => temp(5549 DOWNTO 5540) := ADC(11 DOWNTO 2);
			WHEN 555 => temp(5559 DOWNTO 5550) := ADC(11 DOWNTO 2);
			WHEN 556 => temp(5569 DOWNTO 5560) := ADC(11 DOWNTO 2);
			WHEN 557 => temp(5579 DOWNTO 5570) := ADC(11 DOWNTO 2);
			WHEN 558 => temp(5589 DOWNTO 5580) := ADC(11 DOWNTO 2);
			WHEN 559 => temp(5599 DOWNTO 5590) := ADC(11 DOWNTO 2);
			WHEN 560 => temp(5609 DOWNTO 5600) := ADC(11 DOWNTO 2);
			WHEN 561 => temp(5619 DOWNTO 5610) := ADC(11 DOWNTO 2);
			WHEN 562 => temp(5629 DOWNTO 5620) := ADC(11 DOWNTO 2);
			WHEN 563 => temp(5639 DOWNTO 5630) := ADC(11 DOWNTO 2);
			WHEN 564 => temp(5649 DOWNTO 5640) := ADC(11 DOWNTO 2);
			WHEN 565 => temp(5659 DOWNTO 5650) := ADC(11 DOWNTO 2);
			WHEN 566 => temp(5669 DOWNTO 5660) := ADC(11 DOWNTO 2);
			WHEN 567 => temp(5679 DOWNTO 5670) := ADC(11 DOWNTO 2);
			WHEN 568 => temp(5689 DOWNTO 5680) := ADC(11 DOWNTO 2);
			WHEN 569 => temp(5699 DOWNTO 5690) := ADC(11 DOWNTO 2);
			WHEN 570 => temp(5709 DOWNTO 5700) := ADC(11 DOWNTO 2);
			WHEN 571 => temp(5719 DOWNTO 5710) := ADC(11 DOWNTO 2);
			WHEN 572 => temp(5729 DOWNTO 5720) := ADC(11 DOWNTO 2);
			WHEN 573 => temp(5739 DOWNTO 5730) := ADC(11 DOWNTO 2);
			WHEN 574 => temp(5749 DOWNTO 5740) := ADC(11 DOWNTO 2);
			WHEN 575 => temp(5759 DOWNTO 5750) := ADC(11 DOWNTO 2);
			WHEN 576 => temp(5769 DOWNTO 5760) := ADC(11 DOWNTO 2);
			WHEN 577 => temp(5779 DOWNTO 5770) := ADC(11 DOWNTO 2);
			WHEN 578 => temp(5789 DOWNTO 5780) := ADC(11 DOWNTO 2);
			WHEN 579 => temp(5799 DOWNTO 5790) := ADC(11 DOWNTO 2);
			WHEN 580 => temp(5809 DOWNTO 5800) := ADC(11 DOWNTO 2);
			WHEN 581 => temp(5819 DOWNTO 5810) := ADC(11 DOWNTO 2);
			WHEN 582 => temp(5829 DOWNTO 5820) := ADC(11 DOWNTO 2);
			WHEN 583 => temp(5839 DOWNTO 5830) := ADC(11 DOWNTO 2);
			WHEN 584 => temp(5849 DOWNTO 5840) := ADC(11 DOWNTO 2);
			WHEN 585 => temp(5859 DOWNTO 5850) := ADC(11 DOWNTO 2);
			WHEN 586 => temp(5869 DOWNTO 5860) := ADC(11 DOWNTO 2);
			WHEN 587 => temp(5879 DOWNTO 5870) := ADC(11 DOWNTO 2);
			WHEN 588 => temp(5889 DOWNTO 5880) := ADC(11 DOWNTO 2);
			WHEN 589 => temp(5899 DOWNTO 5890) := ADC(11 DOWNTO 2);
			WHEN 590 => temp(5909 DOWNTO 5900) := ADC(11 DOWNTO 2);
			WHEN 591 => temp(5919 DOWNTO 5910) := ADC(11 DOWNTO 2);
			WHEN 592 => temp(5929 DOWNTO 5920) := ADC(11 DOWNTO 2);
			WHEN 593 => temp(5939 DOWNTO 5930) := ADC(11 DOWNTO 2);
			WHEN 594 => temp(5949 DOWNTO 5940) := ADC(11 DOWNTO 2);
			WHEN 595 => temp(5959 DOWNTO 5950) := ADC(11 DOWNTO 2);
			WHEN 596 => temp(5969 DOWNTO 5960) := ADC(11 DOWNTO 2);
			WHEN 597 => temp(5979 DOWNTO 5970) := ADC(11 DOWNTO 2);
			WHEN 598 => temp(5989 DOWNTO 5980) := ADC(11 DOWNTO 2);
			WHEN 599 => temp(5999 DOWNTO 5990) := ADC(11 DOWNTO 2);
			WHEN 600 => temp(6009 DOWNTO 6000) := ADC(11 DOWNTO 2);
			WHEN 601 => temp(6019 DOWNTO 6010) := ADC(11 DOWNTO 2);
			WHEN 602 => temp(6029 DOWNTO 6020) := ADC(11 DOWNTO 2);
			WHEN 603 => temp(6039 DOWNTO 6030) := ADC(11 DOWNTO 2);
			WHEN 604 => temp(6049 DOWNTO 6040) := ADC(11 DOWNTO 2);
			WHEN 605 => temp(6059 DOWNTO 6050) := ADC(11 DOWNTO 2);
			WHEN 606 => temp(6069 DOWNTO 6060) := ADC(11 DOWNTO 2);
			WHEN 607 => temp(6079 DOWNTO 6070) := ADC(11 DOWNTO 2);
			WHEN 608 => temp(6089 DOWNTO 6080) := ADC(11 DOWNTO 2);
			WHEN 609 => temp(6099 DOWNTO 6090) := ADC(11 DOWNTO 2);
			WHEN 610 => temp(6109 DOWNTO 6100) := ADC(11 DOWNTO 2);
			WHEN 611 => temp(6119 DOWNTO 6110) := ADC(11 DOWNTO 2);
			WHEN 612 => temp(6129 DOWNTO 6120) := ADC(11 DOWNTO 2);
			WHEN 613 => temp(6139 DOWNTO 6130) := ADC(11 DOWNTO 2);
			WHEN 614 => temp(6149 DOWNTO 6140) := ADC(11 DOWNTO 2);
			WHEN 615 => temp(6159 DOWNTO 6150) := ADC(11 DOWNTO 2);
			WHEN 616 => temp(6169 DOWNTO 6160) := ADC(11 DOWNTO 2);
			WHEN 617 => temp(6179 DOWNTO 6170) := ADC(11 DOWNTO 2);
			WHEN 618 => temp(6189 DOWNTO 6180) := ADC(11 DOWNTO 2);
			WHEN 619 => temp(6199 DOWNTO 6190) := ADC(11 DOWNTO 2);
			WHEN 620 => temp(6209 DOWNTO 6200) := ADC(11 DOWNTO 2);
			WHEN 621 => temp(6219 DOWNTO 6210) := ADC(11 DOWNTO 2);
			WHEN 622 => temp(6229 DOWNTO 6220) := ADC(11 DOWNTO 2);
			WHEN 623 => temp(6239 DOWNTO 6230) := ADC(11 DOWNTO 2);
			WHEN 624 => temp(6249 DOWNTO 6240) := ADC(11 DOWNTO 2);
			WHEN 625 => temp(6259 DOWNTO 6250) := ADC(11 DOWNTO 2);
			WHEN 626 => temp(6269 DOWNTO 6260) := ADC(11 DOWNTO 2);
			WHEN 627 => temp(6279 DOWNTO 6270) := ADC(11 DOWNTO 2);
			WHEN 628 => temp(6289 DOWNTO 6280) := ADC(11 DOWNTO 2);
			WHEN 629 => temp(6299 DOWNTO 6290) := ADC(11 DOWNTO 2);
			WHEN 630 => temp(6309 DOWNTO 6300) := ADC(11 DOWNTO 2);
			WHEN 631 => temp(6319 DOWNTO 6310) := ADC(11 DOWNTO 2);
			WHEN 632 => temp(6329 DOWNTO 6320) := ADC(11 DOWNTO 2);
			WHEN 633 => temp(6339 DOWNTO 6330) := ADC(11 DOWNTO 2);
			WHEN 634 => temp(6349 DOWNTO 6340) := ADC(11 DOWNTO 2);
			WHEN 635 => temp(6359 DOWNTO 6350) := ADC(11 DOWNTO 2);
			WHEN 636 => temp(6369 DOWNTO 6360) := ADC(11 DOWNTO 2);
			WHEN 637 => temp(6379 DOWNTO 6370) := ADC(11 DOWNTO 2);
			WHEN 638 => temp(6389 DOWNTO 6380) := ADC(11 DOWNTO 2);
			WHEN 639 => temp(6399 DOWNTO 6390) := ADC(11 DOWNTO 2);
			WHEN 640 => temp(6409 DOWNTO 6400) := ADC(11 DOWNTO 2);
			WHEN 641 => temp(6419 DOWNTO 6410) := ADC(11 DOWNTO 2);
			WHEN 642 => temp(6429 DOWNTO 6420) := ADC(11 DOWNTO 2);
			WHEN 643 => temp(6439 DOWNTO 6430) := ADC(11 DOWNTO 2);
			WHEN 644 => temp(6449 DOWNTO 6440) := ADC(11 DOWNTO 2);
			WHEN 645 => temp(6459 DOWNTO 6450) := ADC(11 DOWNTO 2);
			WHEN 646 => temp(6469 DOWNTO 6460) := ADC(11 DOWNTO 2);
			WHEN 647 => temp(6479 DOWNTO 6470) := ADC(11 DOWNTO 2);
			WHEN 648 => temp(6489 DOWNTO 6480) := ADC(11 DOWNTO 2);
			WHEN 649 => temp(6499 DOWNTO 6490) := ADC(11 DOWNTO 2);
			WHEN 650 => temp(6509 DOWNTO 6500) := ADC(11 DOWNTO 2);
			WHEN 651 => temp(6519 DOWNTO 6510) := ADC(11 DOWNTO 2);
			WHEN 652 => temp(6529 DOWNTO 6520) := ADC(11 DOWNTO 2);
			WHEN 653 => temp(6539 DOWNTO 6530) := ADC(11 DOWNTO 2);
			WHEN 654 => temp(6549 DOWNTO 6540) := ADC(11 DOWNTO 2);
			WHEN 655 => temp(6559 DOWNTO 6550) := ADC(11 DOWNTO 2);
			WHEN 656 => temp(6569 DOWNTO 6560) := ADC(11 DOWNTO 2);
			WHEN 657 => temp(6579 DOWNTO 6570) := ADC(11 DOWNTO 2);
			WHEN 658 => temp(6589 DOWNTO 6580) := ADC(11 DOWNTO 2);
			WHEN 659 => temp(6599 DOWNTO 6590) := ADC(11 DOWNTO 2);
			WHEN 660 => temp(6609 DOWNTO 6600) := ADC(11 DOWNTO 2);
			WHEN 661 => temp(6619 DOWNTO 6610) := ADC(11 DOWNTO 2);
			WHEN 662 => temp(6629 DOWNTO 6620) := ADC(11 DOWNTO 2);
			WHEN 663 => temp(6639 DOWNTO 6630) := ADC(11 DOWNTO 2);
			WHEN 664 => temp(6649 DOWNTO 6640) := ADC(11 DOWNTO 2);
			WHEN 665 => temp(6659 DOWNTO 6650) := ADC(11 DOWNTO 2);
			WHEN 666 => temp(6669 DOWNTO 6660) := ADC(11 DOWNTO 2);
			WHEN 667 => temp(6679 DOWNTO 6670) := ADC(11 DOWNTO 2);
			WHEN 668 => temp(6689 DOWNTO 6680) := ADC(11 DOWNTO 2);
			WHEN 669 => temp(6699 DOWNTO 6690) := ADC(11 DOWNTO 2);
			WHEN 670 => temp(6709 DOWNTO 6700) := ADC(11 DOWNTO 2);
			WHEN 671 => temp(6719 DOWNTO 6710) := ADC(11 DOWNTO 2);
			WHEN 672 => temp(6729 DOWNTO 6720) := ADC(11 DOWNTO 2);
			WHEN 673 => temp(6739 DOWNTO 6730) := ADC(11 DOWNTO 2);
			WHEN 674 => temp(6749 DOWNTO 6740) := ADC(11 DOWNTO 2);
			WHEN 675 => temp(6759 DOWNTO 6750) := ADC(11 DOWNTO 2);
			WHEN 676 => temp(6769 DOWNTO 6760) := ADC(11 DOWNTO 2);
			WHEN 677 => temp(6779 DOWNTO 6770) := ADC(11 DOWNTO 2);
			WHEN 678 => temp(6789 DOWNTO 6780) := ADC(11 DOWNTO 2);
			WHEN 679 => temp(6799 DOWNTO 6790) := ADC(11 DOWNTO 2);
			WHEN 680 => temp(6809 DOWNTO 6800) := ADC(11 DOWNTO 2);
			WHEN 681 => temp(6819 DOWNTO 6810) := ADC(11 DOWNTO 2);
			WHEN 682 => temp(6829 DOWNTO 6820) := ADC(11 DOWNTO 2);
			WHEN 683 => temp(6839 DOWNTO 6830) := ADC(11 DOWNTO 2);
			WHEN 684 => temp(6849 DOWNTO 6840) := ADC(11 DOWNTO 2);
			WHEN 685 => temp(6859 DOWNTO 6850) := ADC(11 DOWNTO 2);
			WHEN 686 => temp(6869 DOWNTO 6860) := ADC(11 DOWNTO 2);
			WHEN 687 => temp(6879 DOWNTO 6870) := ADC(11 DOWNTO 2);
			WHEN 688 => temp(6889 DOWNTO 6880) := ADC(11 DOWNTO 2);
			WHEN 689 => temp(6899 DOWNTO 6890) := ADC(11 DOWNTO 2);
			WHEN 690 => temp(6909 DOWNTO 6900) := ADC(11 DOWNTO 2);
			WHEN 691 => temp(6919 DOWNTO 6910) := ADC(11 DOWNTO 2);
			WHEN 692 => temp(6929 DOWNTO 6920) := ADC(11 DOWNTO 2);
			WHEN 693 => temp(6939 DOWNTO 6930) := ADC(11 DOWNTO 2);
			WHEN 694 => temp(6949 DOWNTO 6940) := ADC(11 DOWNTO 2);
			WHEN 695 => temp(6959 DOWNTO 6950) := ADC(11 DOWNTO 2);
			WHEN 696 => temp(6969 DOWNTO 6960) := ADC(11 DOWNTO 2);
			WHEN 697 => temp(6979 DOWNTO 6970) := ADC(11 DOWNTO 2);
			WHEN 698 => temp(6989 DOWNTO 6980) := ADC(11 DOWNTO 2);
			WHEN 699 => temp(6999 DOWNTO 6990) := ADC(11 DOWNTO 2);
			WHEN 700 => temp(7009 DOWNTO 7000) := ADC(11 DOWNTO 2);
			WHEN 701 => temp(7019 DOWNTO 7010) := ADC(11 DOWNTO 2);
			WHEN 702 => temp(7029 DOWNTO 7020) := ADC(11 DOWNTO 2);
			WHEN 703 => temp(7039 DOWNTO 7030) := ADC(11 DOWNTO 2);
			WHEN 704 => temp(7049 DOWNTO 7040) := ADC(11 DOWNTO 2);
			WHEN 705 => temp(7059 DOWNTO 7050) := ADC(11 DOWNTO 2);
			WHEN 706 => temp(7069 DOWNTO 7060) := ADC(11 DOWNTO 2);
			WHEN 707 => temp(7079 DOWNTO 7070) := ADC(11 DOWNTO 2);
			WHEN 708 => temp(7089 DOWNTO 7080) := ADC(11 DOWNTO 2);
			WHEN 709 => temp(7099 DOWNTO 7090) := ADC(11 DOWNTO 2);
			WHEN 710 => temp(7109 DOWNTO 7100) := ADC(11 DOWNTO 2);
			WHEN 711 => temp(7119 DOWNTO 7110) := ADC(11 DOWNTO 2);
			WHEN 712 => temp(7129 DOWNTO 7120) := ADC(11 DOWNTO 2);
			WHEN 713 => temp(7139 DOWNTO 7130) := ADC(11 DOWNTO 2);
			WHEN 714 => temp(7149 DOWNTO 7140) := ADC(11 DOWNTO 2);
			WHEN 715 => temp(7159 DOWNTO 7150) := ADC(11 DOWNTO 2);
			WHEN 716 => temp(7169 DOWNTO 7160) := ADC(11 DOWNTO 2);
			WHEN 717 => temp(7179 DOWNTO 7170) := ADC(11 DOWNTO 2);
			WHEN 718 => temp(7189 DOWNTO 7180) := ADC(11 DOWNTO 2);
			WHEN 719 => temp(7199 DOWNTO 7190) := ADC(11 DOWNTO 2);
			WHEN 720 => temp(7209 DOWNTO 7200) := ADC(11 DOWNTO 2);
			WHEN 721 => temp(7219 DOWNTO 7210) := ADC(11 DOWNTO 2);
			WHEN 722 => temp(7229 DOWNTO 7220) := ADC(11 DOWNTO 2);
			WHEN 723 => temp(7239 DOWNTO 7230) := ADC(11 DOWNTO 2);
			WHEN 724 => temp(7249 DOWNTO 7240) := ADC(11 DOWNTO 2);
			WHEN 725 => temp(7259 DOWNTO 7250) := ADC(11 DOWNTO 2);
			WHEN 726 => temp(7269 DOWNTO 7260) := ADC(11 DOWNTO 2);
			WHEN 727 => temp(7279 DOWNTO 7270) := ADC(11 DOWNTO 2);
			WHEN 728 => temp(7289 DOWNTO 7280) := ADC(11 DOWNTO 2);
			WHEN 729 => temp(7299 DOWNTO 7290) := ADC(11 DOWNTO 2);
			WHEN 730 => temp(7309 DOWNTO 7300) := ADC(11 DOWNTO 2);
			WHEN 731 => temp(7319 DOWNTO 7310) := ADC(11 DOWNTO 2);
			WHEN 732 => temp(7329 DOWNTO 7320) := ADC(11 DOWNTO 2);
			WHEN 733 => temp(7339 DOWNTO 7330) := ADC(11 DOWNTO 2);
			WHEN 734 => temp(7349 DOWNTO 7340) := ADC(11 DOWNTO 2);
			WHEN 735 => temp(7359 DOWNTO 7350) := ADC(11 DOWNTO 2);
			WHEN 736 => temp(7369 DOWNTO 7360) := ADC(11 DOWNTO 2);
			WHEN 737 => temp(7379 DOWNTO 7370) := ADC(11 DOWNTO 2);
			WHEN 738 => temp(7389 DOWNTO 7380) := ADC(11 DOWNTO 2);
			WHEN 739 => temp(7399 DOWNTO 7390) := ADC(11 DOWNTO 2);
			WHEN 740 => temp(7409 DOWNTO 7400) := ADC(11 DOWNTO 2);
			WHEN 741 => temp(7419 DOWNTO 7410) := ADC(11 DOWNTO 2);
			WHEN 742 => temp(7429 DOWNTO 7420) := ADC(11 DOWNTO 2);
			WHEN 743 => temp(7439 DOWNTO 7430) := ADC(11 DOWNTO 2);
			WHEN 744 => temp(7449 DOWNTO 7440) := ADC(11 DOWNTO 2);
			WHEN 745 => temp(7459 DOWNTO 7450) := ADC(11 DOWNTO 2);
			WHEN 746 => temp(7469 DOWNTO 7460) := ADC(11 DOWNTO 2);
			WHEN 747 => temp(7479 DOWNTO 7470) := ADC(11 DOWNTO 2);
			WHEN 748 => temp(7489 DOWNTO 7480) := ADC(11 DOWNTO 2);
			WHEN 749 => temp(7499 DOWNTO 7490) := ADC(11 DOWNTO 2);
			WHEN 750 => temp(7509 DOWNTO 7500) := ADC(11 DOWNTO 2);
			WHEN 751 => temp(7519 DOWNTO 7510) := ADC(11 DOWNTO 2);
			WHEN 752 => temp(7529 DOWNTO 7520) := ADC(11 DOWNTO 2);
			WHEN 753 => temp(7539 DOWNTO 7530) := ADC(11 DOWNTO 2);
			WHEN 754 => temp(7549 DOWNTO 7540) := ADC(11 DOWNTO 2);
			WHEN 755 => temp(7559 DOWNTO 7550) := ADC(11 DOWNTO 2);
			WHEN 756 => temp(7569 DOWNTO 7560) := ADC(11 DOWNTO 2);
			WHEN 757 => temp(7579 DOWNTO 7570) := ADC(11 DOWNTO 2);
			WHEN 758 => temp(7589 DOWNTO 7580) := ADC(11 DOWNTO 2);
			WHEN 759 => temp(7599 DOWNTO 7590) := ADC(11 DOWNTO 2);
			WHEN 760 => temp(7609 DOWNTO 7600) := ADC(11 DOWNTO 2);
			WHEN 761 => temp(7619 DOWNTO 7610) := ADC(11 DOWNTO 2);
			WHEN 762 => temp(7629 DOWNTO 7620) := ADC(11 DOWNTO 2);
			WHEN 763 => temp(7639 DOWNTO 7630) := ADC(11 DOWNTO 2);
			WHEN 764 => temp(7649 DOWNTO 7640) := ADC(11 DOWNTO 2);
			WHEN 765 => temp(7659 DOWNTO 7650) := ADC(11 DOWNTO 2);
			WHEN 766 => temp(7669 DOWNTO 7660) := ADC(11 DOWNTO 2);
			WHEN 767 => temp(7679 DOWNTO 7670) := ADC(11 DOWNTO 2);
			WHEN 768 => temp(7689 DOWNTO 7680) := ADC(11 DOWNTO 2);
			WHEN 769 => temp(7699 DOWNTO 7690) := ADC(11 DOWNTO 2);
			WHEN 770 => temp(7709 DOWNTO 7700) := ADC(11 DOWNTO 2);
			WHEN 771 => temp(7719 DOWNTO 7710) := ADC(11 DOWNTO 2);
			WHEN 772 => temp(7729 DOWNTO 7720) := ADC(11 DOWNTO 2);
			WHEN 773 => temp(7739 DOWNTO 7730) := ADC(11 DOWNTO 2);
			WHEN 774 => temp(7749 DOWNTO 7740) := ADC(11 DOWNTO 2);
			WHEN 775 => temp(7759 DOWNTO 7750) := ADC(11 DOWNTO 2);
			WHEN 776 => temp(7769 DOWNTO 7760) := ADC(11 DOWNTO 2);
			WHEN 777 => temp(7779 DOWNTO 7770) := ADC(11 DOWNTO 2);
			WHEN 778 => temp(7789 DOWNTO 7780) := ADC(11 DOWNTO 2);
			WHEN 779 => temp(7799 DOWNTO 7790) := ADC(11 DOWNTO 2);
			WHEN 780 => temp(7809 DOWNTO 7800) := ADC(11 DOWNTO 2);
			WHEN 781 => temp(7819 DOWNTO 7810) := ADC(11 DOWNTO 2);
			WHEN 782 => temp(7829 DOWNTO 7820) := ADC(11 DOWNTO 2);
			WHEN 783 => temp(7839 DOWNTO 7830) := ADC(11 DOWNTO 2);
			WHEN 784 => temp(7849 DOWNTO 7840) := ADC(11 DOWNTO 2);
			WHEN 785 => temp(7859 DOWNTO 7850) := ADC(11 DOWNTO 2);
			WHEN 786 => temp(7869 DOWNTO 7860) := ADC(11 DOWNTO 2);
			WHEN 787 => temp(7879 DOWNTO 7870) := ADC(11 DOWNTO 2);
			WHEN 788 => temp(7889 DOWNTO 7880) := ADC(11 DOWNTO 2);
			WHEN 789 => temp(7899 DOWNTO 7890) := ADC(11 DOWNTO 2);
			WHEN 790 => temp(7909 DOWNTO 7900) := ADC(11 DOWNTO 2);
			WHEN 791 => temp(7919 DOWNTO 7910) := ADC(11 DOWNTO 2);
			WHEN 792 => temp(7929 DOWNTO 7920) := ADC(11 DOWNTO 2);
			WHEN 793 => temp(7939 DOWNTO 7930) := ADC(11 DOWNTO 2);
			WHEN 794 => temp(7949 DOWNTO 7940) := ADC(11 DOWNTO 2);
			WHEN 795 => temp(7959 DOWNTO 7950) := ADC(11 DOWNTO 2);
			WHEN 796 => temp(7969 DOWNTO 7960) := ADC(11 DOWNTO 2);
			WHEN 797 => temp(7979 DOWNTO 7970) := ADC(11 DOWNTO 2);
			WHEN 798 => temp(7989 DOWNTO 7980) := ADC(11 DOWNTO 2);
			WHEN 799 => temp(7999 DOWNTO 7990) := ADC(11 DOWNTO 2);
			WHEN 800 => temp(8009 DOWNTO 8000) := ADC(11 DOWNTO 2);
			WHEN 801 => temp(8019 DOWNTO 8010) := ADC(11 DOWNTO 2);
			WHEN 802 => temp(8029 DOWNTO 8020) := ADC(11 DOWNTO 2);
			WHEN 803 => temp(8039 DOWNTO 8030) := ADC(11 DOWNTO 2);
			WHEN 804 => temp(8049 DOWNTO 8040) := ADC(11 DOWNTO 2);
			WHEN 805 => temp(8059 DOWNTO 8050) := ADC(11 DOWNTO 2);
			WHEN 806 => temp(8069 DOWNTO 8060) := ADC(11 DOWNTO 2);
			WHEN 807 => temp(8079 DOWNTO 8070) := ADC(11 DOWNTO 2);
			WHEN 808 => temp(8089 DOWNTO 8080) := ADC(11 DOWNTO 2);
			WHEN 809 => temp(8099 DOWNTO 8090) := ADC(11 DOWNTO 2);
			WHEN 810 => temp(8109 DOWNTO 8100) := ADC(11 DOWNTO 2);
			WHEN 811 => temp(8119 DOWNTO 8110) := ADC(11 DOWNTO 2);
			WHEN 812 => temp(8129 DOWNTO 8120) := ADC(11 DOWNTO 2);
			WHEN 813 => temp(8139 DOWNTO 8130) := ADC(11 DOWNTO 2);
			WHEN 814 => temp(8149 DOWNTO 8140) := ADC(11 DOWNTO 2);
			WHEN 815 => temp(8159 DOWNTO 8150) := ADC(11 DOWNTO 2);
			WHEN 816 => temp(8169 DOWNTO 8160) := ADC(11 DOWNTO 2);
			WHEN 817 => temp(8179 DOWNTO 8170) := ADC(11 DOWNTO 2);
			WHEN 818 => temp(8189 DOWNTO 8180) := ADC(11 DOWNTO 2);
			WHEN 819 => temp(8199 DOWNTO 8190) := ADC(11 DOWNTO 2);
			WHEN 820 => temp(8209 DOWNTO 8200) := ADC(11 DOWNTO 2);
			WHEN 821 => temp(8219 DOWNTO 8210) := ADC(11 DOWNTO 2);
			WHEN 822 => temp(8229 DOWNTO 8220) := ADC(11 DOWNTO 2);
			WHEN 823 => temp(8239 DOWNTO 8230) := ADC(11 DOWNTO 2);
			WHEN 824 => temp(8249 DOWNTO 8240) := ADC(11 DOWNTO 2);
			WHEN 825 => temp(8259 DOWNTO 8250) := ADC(11 DOWNTO 2);
			WHEN 826 => temp(8269 DOWNTO 8260) := ADC(11 DOWNTO 2);
			WHEN 827 => temp(8279 DOWNTO 8270) := ADC(11 DOWNTO 2);
			WHEN 828 => temp(8289 DOWNTO 8280) := ADC(11 DOWNTO 2);
			WHEN 829 => temp(8299 DOWNTO 8290) := ADC(11 DOWNTO 2);
			WHEN 830 => temp(8309 DOWNTO 8300) := ADC(11 DOWNTO 2);
			WHEN 831 => temp(8319 DOWNTO 8310) := ADC(11 DOWNTO 2);
			WHEN 832 => temp(8329 DOWNTO 8320) := ADC(11 DOWNTO 2);
			WHEN 833 => temp(8339 DOWNTO 8330) := ADC(11 DOWNTO 2);
			WHEN 834 => temp(8349 DOWNTO 8340) := ADC(11 DOWNTO 2);
			WHEN 835 => temp(8359 DOWNTO 8350) := ADC(11 DOWNTO 2);
			WHEN 836 => temp(8369 DOWNTO 8360) := ADC(11 DOWNTO 2);
			WHEN 837 => temp(8379 DOWNTO 8370) := ADC(11 DOWNTO 2);
			WHEN 838 => temp(8389 DOWNTO 8380) := ADC(11 DOWNTO 2);
			WHEN 839 => temp(8399 DOWNTO 8390) := ADC(11 DOWNTO 2);
			WHEN 840 => temp(8409 DOWNTO 8400) := ADC(11 DOWNTO 2);
			WHEN 841 => temp(8419 DOWNTO 8410) := ADC(11 DOWNTO 2);
			WHEN 842 => temp(8429 DOWNTO 8420) := ADC(11 DOWNTO 2);
			WHEN 843 => temp(8439 DOWNTO 8430) := ADC(11 DOWNTO 2);
			WHEN 844 => temp(8449 DOWNTO 8440) := ADC(11 DOWNTO 2);
			WHEN 845 => temp(8459 DOWNTO 8450) := ADC(11 DOWNTO 2);
			WHEN 846 => temp(8469 DOWNTO 8460) := ADC(11 DOWNTO 2);
			WHEN 847 => temp(8479 DOWNTO 8470) := ADC(11 DOWNTO 2);
			WHEN 848 => temp(8489 DOWNTO 8480) := ADC(11 DOWNTO 2);
			WHEN 849 => temp(8499 DOWNTO 8490) := ADC(11 DOWNTO 2);
			WHEN 850 => temp(8509 DOWNTO 8500) := ADC(11 DOWNTO 2);
			WHEN 851 => temp(8519 DOWNTO 8510) := ADC(11 DOWNTO 2);
			WHEN 852 => temp(8529 DOWNTO 8520) := ADC(11 DOWNTO 2);
			WHEN 853 => temp(8539 DOWNTO 8530) := ADC(11 DOWNTO 2);
			WHEN 854 => temp(8549 DOWNTO 8540) := ADC(11 DOWNTO 2);
			WHEN 855 => temp(8559 DOWNTO 8550) := ADC(11 DOWNTO 2);
			WHEN 856 => temp(8569 DOWNTO 8560) := ADC(11 DOWNTO 2);
			WHEN 857 => temp(8579 DOWNTO 8570) := ADC(11 DOWNTO 2);
			WHEN 858 => temp(8589 DOWNTO 8580) := ADC(11 DOWNTO 2);
			WHEN 859 => temp(8599 DOWNTO 8590) := ADC(11 DOWNTO 2);
			WHEN 860 => temp(8609 DOWNTO 8600) := ADC(11 DOWNTO 2);
			WHEN 861 => temp(8619 DOWNTO 8610) := ADC(11 DOWNTO 2);
			WHEN 862 => temp(8629 DOWNTO 8620) := ADC(11 DOWNTO 2);
			WHEN 863 => temp(8639 DOWNTO 8630) := ADC(11 DOWNTO 2);
			WHEN 864 => temp(8649 DOWNTO 8640) := ADC(11 DOWNTO 2);
			WHEN 865 => temp(8659 DOWNTO 8650) := ADC(11 DOWNTO 2);
			WHEN 866 => temp(8669 DOWNTO 8660) := ADC(11 DOWNTO 2);
			WHEN 867 => temp(8679 DOWNTO 8670) := ADC(11 DOWNTO 2);
			WHEN 868 => temp(8689 DOWNTO 8680) := ADC(11 DOWNTO 2);
			WHEN 869 => temp(8699 DOWNTO 8690) := ADC(11 DOWNTO 2);
			WHEN 870 => temp(8709 DOWNTO 8700) := ADC(11 DOWNTO 2);
			WHEN 871 => temp(8719 DOWNTO 8710) := ADC(11 DOWNTO 2);
			WHEN 872 => temp(8729 DOWNTO 8720) := ADC(11 DOWNTO 2);
			WHEN 873 => temp(8739 DOWNTO 8730) := ADC(11 DOWNTO 2);
			WHEN 874 => temp(8749 DOWNTO 8740) := ADC(11 DOWNTO 2);
			WHEN 875 => temp(8759 DOWNTO 8750) := ADC(11 DOWNTO 2);
			WHEN 876 => temp(8769 DOWNTO 8760) := ADC(11 DOWNTO 2);
			WHEN 877 => temp(8779 DOWNTO 8770) := ADC(11 DOWNTO 2);
			WHEN 878 => temp(8789 DOWNTO 8780) := ADC(11 DOWNTO 2);
			WHEN 879 => temp(8799 DOWNTO 8790) := ADC(11 DOWNTO 2);
			WHEN 880 => temp(8809 DOWNTO 8800) := ADC(11 DOWNTO 2);
			WHEN 881 => temp(8819 DOWNTO 8810) := ADC(11 DOWNTO 2);
			WHEN 882 => temp(8829 DOWNTO 8820) := ADC(11 DOWNTO 2);
			WHEN 883 => temp(8839 DOWNTO 8830) := ADC(11 DOWNTO 2);
			WHEN 884 => temp(8849 DOWNTO 8840) := ADC(11 DOWNTO 2);
			WHEN 885 => temp(8859 DOWNTO 8850) := ADC(11 DOWNTO 2);
			WHEN 886 => temp(8869 DOWNTO 8860) := ADC(11 DOWNTO 2);
			WHEN 887 => temp(8879 DOWNTO 8870) := ADC(11 DOWNTO 2);
			WHEN 888 => temp(8889 DOWNTO 8880) := ADC(11 DOWNTO 2);
			WHEN 889 => temp(8899 DOWNTO 8890) := ADC(11 DOWNTO 2);
			WHEN 890 => temp(8909 DOWNTO 8900) := ADC(11 DOWNTO 2);
			WHEN 891 => temp(8919 DOWNTO 8910) := ADC(11 DOWNTO 2);
			WHEN 892 => temp(8929 DOWNTO 8920) := ADC(11 DOWNTO 2);
			WHEN 893 => temp(8939 DOWNTO 8930) := ADC(11 DOWNTO 2);
			WHEN 894 => temp(8949 DOWNTO 8940) := ADC(11 DOWNTO 2);
			WHEN 895 => temp(8959 DOWNTO 8950) := ADC(11 DOWNTO 2);
			WHEN 896 => temp(8969 DOWNTO 8960) := ADC(11 DOWNTO 2);
			WHEN 897 => temp(8979 DOWNTO 8970) := ADC(11 DOWNTO 2);
			WHEN 898 => temp(8989 DOWNTO 8980) := ADC(11 DOWNTO 2);
			WHEN 899 => temp(8999 DOWNTO 8990) := ADC(11 DOWNTO 2);
			WHEN 900 => temp(9009 DOWNTO 9000) := ADC(11 DOWNTO 2);
			WHEN 901 => temp(9019 DOWNTO 9010) := ADC(11 DOWNTO 2);
			WHEN 902 => temp(9029 DOWNTO 9020) := ADC(11 DOWNTO 2);
			WHEN 903 => temp(9039 DOWNTO 9030) := ADC(11 DOWNTO 2);
			WHEN 904 => temp(9049 DOWNTO 9040) := ADC(11 DOWNTO 2);
			WHEN 905 => temp(9059 DOWNTO 9050) := ADC(11 DOWNTO 2);
			WHEN 906 => temp(9069 DOWNTO 9060) := ADC(11 DOWNTO 2);
			WHEN 907 => temp(9079 DOWNTO 9070) := ADC(11 DOWNTO 2);
			WHEN 908 => temp(9089 DOWNTO 9080) := ADC(11 DOWNTO 2);
			WHEN 909 => temp(9099 DOWNTO 9090) := ADC(11 DOWNTO 2);
			WHEN 910 => temp(9109 DOWNTO 9100) := ADC(11 DOWNTO 2);
			WHEN 911 => temp(9119 DOWNTO 9110) := ADC(11 DOWNTO 2);
			WHEN 912 => temp(9129 DOWNTO 9120) := ADC(11 DOWNTO 2);
			WHEN 913 => temp(9139 DOWNTO 9130) := ADC(11 DOWNTO 2);
			WHEN 914 => temp(9149 DOWNTO 9140) := ADC(11 DOWNTO 2);
			WHEN 915 => temp(9159 DOWNTO 9150) := ADC(11 DOWNTO 2);
			WHEN 916 => temp(9169 DOWNTO 9160) := ADC(11 DOWNTO 2);
			WHEN 917 => temp(9179 DOWNTO 9170) := ADC(11 DOWNTO 2);
			WHEN 918 => temp(9189 DOWNTO 9180) := ADC(11 DOWNTO 2);
			WHEN 919 => temp(9199 DOWNTO 9190) := ADC(11 DOWNTO 2);
			WHEN 920 => temp(9209 DOWNTO 9200) := ADC(11 DOWNTO 2);
			WHEN 921 => temp(9219 DOWNTO 9210) := ADC(11 DOWNTO 2);
			WHEN 922 => temp(9229 DOWNTO 9220) := ADC(11 DOWNTO 2);
			WHEN 923 => temp(9239 DOWNTO 9230) := ADC(11 DOWNTO 2);
			WHEN 924 => temp(9249 DOWNTO 9240) := ADC(11 DOWNTO 2);
			WHEN 925 => temp(9259 DOWNTO 9250) := ADC(11 DOWNTO 2);
			WHEN 926 => temp(9269 DOWNTO 9260) := ADC(11 DOWNTO 2);
			WHEN 927 => temp(9279 DOWNTO 9270) := ADC(11 DOWNTO 2);
			WHEN 928 => temp(9289 DOWNTO 9280) := ADC(11 DOWNTO 2);
			WHEN 929 => temp(9299 DOWNTO 9290) := ADC(11 DOWNTO 2);
			WHEN 930 => temp(9309 DOWNTO 9300) := ADC(11 DOWNTO 2);
			WHEN 931 => temp(9319 DOWNTO 9310) := ADC(11 DOWNTO 2);
			WHEN 932 => temp(9329 DOWNTO 9320) := ADC(11 DOWNTO 2);
			WHEN 933 => temp(9339 DOWNTO 9330) := ADC(11 DOWNTO 2);
			WHEN 934 => temp(9349 DOWNTO 9340) := ADC(11 DOWNTO 2);
			WHEN 935 => temp(9359 DOWNTO 9350) := ADC(11 DOWNTO 2);
			WHEN 936 => temp(9369 DOWNTO 9360) := ADC(11 DOWNTO 2);
			WHEN 937 => temp(9379 DOWNTO 9370) := ADC(11 DOWNTO 2);
			WHEN 938 => temp(9389 DOWNTO 9380) := ADC(11 DOWNTO 2);
			WHEN 939 => temp(9399 DOWNTO 9390) := ADC(11 DOWNTO 2);
			WHEN 940 => temp(9409 DOWNTO 9400) := ADC(11 DOWNTO 2);
			WHEN 941 => temp(9419 DOWNTO 9410) := ADC(11 DOWNTO 2);
			WHEN 942 => temp(9429 DOWNTO 9420) := ADC(11 DOWNTO 2);
			WHEN 943 => temp(9439 DOWNTO 9430) := ADC(11 DOWNTO 2);
			WHEN 944 => temp(9449 DOWNTO 9440) := ADC(11 DOWNTO 2);
			WHEN 945 => temp(9459 DOWNTO 9450) := ADC(11 DOWNTO 2);
			WHEN 946 => temp(9469 DOWNTO 9460) := ADC(11 DOWNTO 2);
			WHEN 947 => temp(9479 DOWNTO 9470) := ADC(11 DOWNTO 2);
			WHEN 948 => temp(9489 DOWNTO 9480) := ADC(11 DOWNTO 2);
			WHEN 949 => temp(9499 DOWNTO 9490) := ADC(11 DOWNTO 2);
			WHEN 950 => temp(9509 DOWNTO 9500) := ADC(11 DOWNTO 2);
			WHEN 951 => temp(9519 DOWNTO 9510) := ADC(11 DOWNTO 2);
			WHEN 952 => temp(9529 DOWNTO 9520) := ADC(11 DOWNTO 2);
			WHEN 953 => temp(9539 DOWNTO 9530) := ADC(11 DOWNTO 2);
			WHEN 954 => temp(9549 DOWNTO 9540) := ADC(11 DOWNTO 2);
			WHEN 955 => temp(9559 DOWNTO 9550) := ADC(11 DOWNTO 2);
			WHEN 956 => temp(9569 DOWNTO 9560) := ADC(11 DOWNTO 2);
			WHEN 957 => temp(9579 DOWNTO 9570) := ADC(11 DOWNTO 2);
			WHEN 958 => temp(9589 DOWNTO 9580) := ADC(11 DOWNTO 2);
			WHEN 959 => temp(9599 DOWNTO 9590) := ADC(11 DOWNTO 2);
			WHEN 960 => temp(9609 DOWNTO 9600) := ADC(11 DOWNTO 2);
			WHEN 961 => temp(9619 DOWNTO 9610) := ADC(11 DOWNTO 2);
			WHEN 962 => temp(9629 DOWNTO 9620) := ADC(11 DOWNTO 2);
			WHEN 963 => temp(9639 DOWNTO 9630) := ADC(11 DOWNTO 2);
			WHEN 964 => temp(9649 DOWNTO 9640) := ADC(11 DOWNTO 2);
			WHEN 965 => temp(9659 DOWNTO 9650) := ADC(11 DOWNTO 2);
			WHEN 966 => temp(9669 DOWNTO 9660) := ADC(11 DOWNTO 2);
			WHEN 967 => temp(9679 DOWNTO 9670) := ADC(11 DOWNTO 2);
			WHEN 968 => temp(9689 DOWNTO 9680) := ADC(11 DOWNTO 2);
			WHEN 969 => temp(9699 DOWNTO 9690) := ADC(11 DOWNTO 2);
			WHEN 970 => temp(9709 DOWNTO 9700) := ADC(11 DOWNTO 2);
			WHEN 971 => temp(9719 DOWNTO 9710) := ADC(11 DOWNTO 2);
			WHEN 972 => temp(9729 DOWNTO 9720) := ADC(11 DOWNTO 2);
			WHEN 973 => temp(9739 DOWNTO 9730) := ADC(11 DOWNTO 2);
			WHEN 974 => temp(9749 DOWNTO 9740) := ADC(11 DOWNTO 2);
			WHEN 975 => temp(9759 DOWNTO 9750) := ADC(11 DOWNTO 2);
			WHEN 976 => temp(9769 DOWNTO 9760) := ADC(11 DOWNTO 2);
			WHEN 977 => temp(9779 DOWNTO 9770) := ADC(11 DOWNTO 2);
			WHEN 978 => temp(9789 DOWNTO 9780) := ADC(11 DOWNTO 2);
			WHEN 979 => temp(9799 DOWNTO 9790) := ADC(11 DOWNTO 2);
			WHEN 980 => temp(9809 DOWNTO 9800) := ADC(11 DOWNTO 2);
			WHEN 981 => temp(9819 DOWNTO 9810) := ADC(11 DOWNTO 2);
			WHEN 982 => temp(9829 DOWNTO 9820) := ADC(11 DOWNTO 2);
			WHEN 983 => temp(9839 DOWNTO 9830) := ADC(11 DOWNTO 2);
			WHEN 984 => temp(9849 DOWNTO 9840) := ADC(11 DOWNTO 2);
			WHEN 985 => temp(9859 DOWNTO 9850) := ADC(11 DOWNTO 2);
			WHEN 986 => temp(9869 DOWNTO 9860) := ADC(11 DOWNTO 2);
			WHEN 987 => temp(9879 DOWNTO 9870) := ADC(11 DOWNTO 2);
			WHEN 988 => temp(9889 DOWNTO 9880) := ADC(11 DOWNTO 2);
			WHEN 989 => temp(9899 DOWNTO 9890) := ADC(11 DOWNTO 2);
			WHEN 990 => temp(9909 DOWNTO 9900) := ADC(11 DOWNTO 2);
			WHEN 991 => temp(9919 DOWNTO 9910) := ADC(11 DOWNTO 2);
			WHEN 992 => temp(9929 DOWNTO 9920) := ADC(11 DOWNTO 2);
			WHEN 993 => temp(9939 DOWNTO 9930) := ADC(11 DOWNTO 2);
			WHEN 994 => temp(9949 DOWNTO 9940) := ADC(11 DOWNTO 2);
			WHEN 995 => temp(9959 DOWNTO 9950) := ADC(11 DOWNTO 2);
			WHEN 996 => temp(9969 DOWNTO 9960) := ADC(11 DOWNTO 2);
			WHEN 997 => temp(9979 DOWNTO 9970) := ADC(11 DOWNTO 2);
			WHEN 998 => temp(9989 DOWNTO 9980) := ADC(11 DOWNTO 2);
			WHEN 999 => temp(9999 DOWNTO 9990) := ADC(11 DOWNTO 2);
			WHEN 1000 => temp(10009 DOWNTO 10000) := ADC(11 DOWNTO 2);
			WHEN 1001 => temp(10019 DOWNTO 10010) := ADC(11 DOWNTO 2);
			WHEN 1002 => temp(10029 DOWNTO 10020) := ADC(11 DOWNTO 2);
			WHEN 1003 => temp(10039 DOWNTO 10030) := ADC(11 DOWNTO 2);
			WHEN 1004 => temp(10049 DOWNTO 10040) := ADC(11 DOWNTO 2);
			WHEN 1005 => temp(10059 DOWNTO 10050) := ADC(11 DOWNTO 2);
			WHEN 1006 => temp(10069 DOWNTO 10060) := ADC(11 DOWNTO 2);
			WHEN 1007 => temp(10079 DOWNTO 10070) := ADC(11 DOWNTO 2);
			WHEN 1008 => temp(10089 DOWNTO 10080) := ADC(11 DOWNTO 2);
			WHEN 1009 => temp(10099 DOWNTO 10090) := ADC(11 DOWNTO 2);
			WHEN 1010 => temp(10109 DOWNTO 10100) := ADC(11 DOWNTO 2);
			WHEN 1011 => temp(10119 DOWNTO 10110) := ADC(11 DOWNTO 2);
			WHEN 1012 => temp(10129 DOWNTO 10120) := ADC(11 DOWNTO 2);
			WHEN 1013 => temp(10139 DOWNTO 10130) := ADC(11 DOWNTO 2);
			WHEN 1014 => temp(10149 DOWNTO 10140) := ADC(11 DOWNTO 2);
			WHEN 1015 => temp(10159 DOWNTO 10150) := ADC(11 DOWNTO 2);
			WHEN 1016 => temp(10169 DOWNTO 10160) := ADC(11 DOWNTO 2);
			WHEN 1017 => temp(10179 DOWNTO 10170) := ADC(11 DOWNTO 2);
			WHEN 1018 => temp(10189 DOWNTO 10180) := ADC(11 DOWNTO 2);
			WHEN 1019 => temp(10199 DOWNTO 10190) := ADC(11 DOWNTO 2);
			WHEN 1020 => temp(10209 DOWNTO 10200) := ADC(11 DOWNTO 2);
			WHEN 1021 => temp(10219 DOWNTO 10210) := ADC(11 DOWNTO 2);
			WHEN 1022 => temp(10229 DOWNTO 10220) := ADC(11 DOWNTO 2);
			WHEN 1023 => temp(10239 DOWNTO 10230) := ADC(11 DOWNTO 2);		
			WHEN OTHERS => NULL;
				END CASE;
			done <= '1';
		ELSE 
			done <= '0';
		END IF;
		samples <= temp;
	END IF;
	END PROCESS;
END;